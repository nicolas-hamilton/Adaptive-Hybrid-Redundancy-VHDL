--| Test31_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:10:10
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test31_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test31_Reg_COMBINED;

architecture a_Test31_Reg_COMBINED of Test31_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 399) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 399) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000");--  398 - 1592

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000011101010000101101", --    2 -    8
      "00000000000000000001010011000011", --    3 -   12
      "00000000000000100001110111000000", --    4 -   16
      "00111000001001000010001100100111", --    5 -   20
      "00000000001001000010100000100101", --    6 -   24
      "00111000010001100000110100110100", --    7 -   28
      "00101100011001110100011001001000", --    8 -   32
      "00100100110010001111010001101010", --    9 -   36
      "00000000110001010100100000000110", --   10 -   40
      "00100001000010101000111000000001", --   11 -   44
      "00000000000001010101100000000111", --   12 -   48
      "00000000110001100110000000000100", --   13 -   52
      "00110101001011010100110100111001", --   14 -   56
      "00000000000011000111000010000011", --   15 -   60
      "10101100000000100000001000111100", --   16 -   64
      "00110001110011110111100111000111", --   17 -   68
      "00000000000000000000000000000000", --   18 -   72
      "00000000000000000000000000000000", --   19 -   76
      "00101001001100001101011001101000", --   20 -   80
      "10101100000001110000001001000000", --   21 -   84
      "00000000000010111000110111000010", --   22 -   88
      "00100110001100101011010101001001", --   23 -   92
      "00000000000000000000000000000000", --   24 -   96
      "00111100000100111000101011001111", --   25 -  100
      "00000000000000000000000000000000", --   26 -  104
      "00000000000100111010010101000010", --   27 -  108
      "00000001101101001010100000100011", --   28 -  112
      "00110100011101100011000000000110", --   29 -  116
      "10101100000010100000001001000100", --   30 -  120
      "00100110000101111111011111011000", --   31 -  124
      "00000000000101111100000110000011", --   32 -  128
      "00000000000000000000000000000000", --   33 -  132
      "10101100000101100000001001001000", --   34 -  136
      "00000010101110001100100000100111", --   35 -  140
      "00000000000000000000000000000000", --   36 -  144
      "10101100000011110000001001001100", --   37 -  148
      "00000010010110011101000000101011", --   38 -  152
      "00000000000000000000000000000000", --   39 -  156
      "10101100000100010000001001010000", --   40 -  160
      "00000000000000000000000000000000", --   41 -  164
      "10101100000110100000001001010100", --   42 -  168
      "00100011111111111111111111111111", --   43 -  172
      "00011111111000001111111111010110", --   44 -  176
      "00010000000000000000000101100001", --   45 -  180
      "00111100000111100000001111100111", --   46 -  184
      "00111100000111110000001111100111", --   47 -  188
      "00000000000111101111010000000010", --   48 -  192
      "00000000000111111111110000000010", --   49 -  196
      "00111100000000011101010000101101", --   50 -  200
      "00111100000011111101010000101101", --   51 -  204
      "00000000000000000001010011000011", --   52 -  208
      "00000000000000001000010011000011", --   53 -  212
      "00000000000000100001110111000000", --   54 -  216
      "00000000000100001000110111000000", --   55 -  220
      "00111000001001000010001100100111", --   56 -  224
      "00111001111100100010001100100111", --   57 -  228
      "00000000001001000010100000100101", --   58 -  232
      "00000001111100101001100000100101", --   59 -  236
      "00111000010001100000110100110100", --   60 -  240
      "00111010000101000000110100110100", --   61 -  244
      "00101100011001110100011001001000", --   62 -  248
      "00101110001101010100011001001000", --   63 -  252
      "00100100110010001111010001101010", --   64 -  256
      "00100110100101101111010001101010", --   65 -  260
      "00000000110001010100100000000110", --   66 -  264
      "00000010100100111011100000000110", --   67 -  268
      "00100001000010101000111000000001", --   68 -  272
      "00100010110110001000111000000001", --   69 -  276
      "00000000000001010101100000000111", --   70 -  280
      "00000000000100111100100000000111", --   71 -  284
      "00000000110001100110000000000100", --   72 -  288
      "00000010100101001101000000000100", --   73 -  292
      "00110101001011010100110100111001", --   74 -  296
      "00110110111110110100110100111001", --   75 -  300
      "00000000000011000111000010000011", --   76 -  304
      "00000000000110101110000010000011", --   77 -  308
      "00010100010100000000000010110011", --   78 -  312
      "10101100000000100000001000111100", --   79 -  316
      "00110001110000010111100111000111", --   80 -  320
      "00110011100011110111100111000111", --   81 -  324
      "00000000000000000000000000000000", --   82 -  328
      "00000000000000000000000000000000", --   83 -  332
      "00000000000000000000000000000000", --   84 -  336
      "00000000000000000000000000000000", --   85 -  340
      "00101001001001001101011001101000", --   86 -  344
      "00101010111100101101011001101000", --   87 -  348
      "00010100111101010000000010101001", --   88 -  352
      "10101100000001110000001001000000", --   89 -  356
      "00000000000010110100010111000010", --   90 -  360
      "00000000000110011011010111000010", --   91 -  364
      "00100101000001011011010101001001", --   92 -  368
      "00100110110100111011010101001001", --   93 -  372
      "00000000000000000000000000000000", --   94 -  376
      "00000000000000000000000000000000", --   95 -  380
      "00111100000001101000101011001111", --   96 -  384
      "00111100000101001000101011001111", --   97 -  388
      "00000000000000000000000000000000", --   98 -  392
      "00000000000000000000000000000000", --   99 -  396
      "00000000000001100110010101000010", --  100 -  400
      "00000000000101001101010101000010", --  101 -  404
      "00000001101011000001000000100011", --  102 -  408
      "00000011011110101000000000100011", --  103 -  412
      "00110100011011100011000000000110", --  104 -  416
      "00110110001111000011000000000110", --  105 -  420
      "00010101010110000000000010010111", --  106 -  424
      "10101100000010100000001001000100", --  107 -  428
      "00100100100010011111011111011000", --  108 -  432
      "00100110010101111111011111011000", --  109 -  436
      "00000000000010010011100110000011", --  110 -  440
      "00000000000101111010100110000011", --  111 -  444
      "00000000000000000000000000000000", --  112 -  448
      "00000000000000000000000000000000", --  113 -  452
      "00010101110111000000000010001111", --  114 -  456
      "10101100000011100000001001001000", --  115 -  460
      "00000000010001110101100000100111", --  116 -  464
      "00000010000101011100100000100111", --  117 -  468
      "00000000000000000000000000000000", --  118 -  472
      "00000000000000000000000000000000", --  119 -  476
      "00010100001011110000000010001001", --  120 -  480
      "10101100000000010000001001001100", --  121 -  484
      "00000000101010110011000000101011", --  122 -  488
      "00000010011110011010000000101011", --  123 -  492
      "00000000000000000000000000000000", --  124 -  496
      "00000000000000000000000000000000", --  125 -  500
      "00010101000101100000000010000011", --  126 -  504
      "10101100000010000000001001010000", --  127 -  508
      "00000000000000000000000000000000", --  128 -  512
      "00000000000000000000000000000000", --  129 -  516
      "00010100110101000000000001111111", --  130 -  520
      "10101100000001100000001001010100", --  131 -  524
      "00100011110111011111111100000110", --  132 -  528
      "00010011101000000000000000010001", --  133 -  532
      "00100011110111011111111000001100", --  134 -  536
      "00010011101000000000000000001111", --  135 -  540
      "00100011110111011111110100010010", --  136 -  544
      "00010011101000000000000000001101", --  137 -  548
      "00100011110111101111111111111111", --  138 -  552
      "00100011111111111111111111111111", --  139 -  556
      "00010111110111110000000001110101", --  140 -  560
      "00011111111000001111111110100101", --  141 -  564
      "00010000000000000000000100000000", --  142 -  568
      "00000000000000000000000000000000", --  143 -  572
      "00000000000000000000000000000000", --  144 -  576
      "00000000000000000000000000000000", --  145 -  580
      "00000000000000000000000000000000", --  146 -  584
      "00000000000000000000000000000000", --  147 -  588
      "00000000000000000000000000000000", --  148 -  592
      "00000000000000000000000000000000", --  149 -  596
      "10001100000111010000010110101100", --  150 -  600
      "00011111101000000000000000000011", --  151 -  604
      "00100000000111010000000000111100", --  152 -  608
      "00010000000000000000000000000010", --  153 -  612
      "00100000000111010000000000000000", --  154 -  616
      "00010100001011110000000001100110", --  155 -  620
      "10101111101000010000010100110100", --  156 -  624
      "10001100000111010000010110101100", --  157 -  628
      "00011111101000000000000000000011", --  158 -  632
      "00100000000111010000000000111100", --  159 -  636
      "00010000000000000000000000000010", --  160 -  640
      "00100000000111010000000000000000", --  161 -  644
      "00010100010100000000000001011111", --  162 -  648
      "10101111101000100000010100111000", --  163 -  652
      "10001100000111010000010110101100", --  164 -  656
      "00011111101000000000000000000011", --  165 -  660
      "00100000000111010000000000111100", --  166 -  664
      "00010000000000000000000000000010", --  167 -  668
      "00100000000111010000000000000000", --  168 -  672
      "00010100011100010000000001011000", --  169 -  676
      "10101111101000110000010100111100", --  170 -  680
      "10001100000111010000010110101100", --  171 -  684
      "00011111101000000000000000000011", --  172 -  688
      "00100000000111010000000000111100", --  173 -  692
      "00010000000000000000000000000010", --  174 -  696
      "00100000000111010000000000000000", --  175 -  700
      "00010100100100100000000001010001", --  176 -  704
      "10101111101001000000010101000000", --  177 -  708
      "10001100000111010000010110101100", --  178 -  712
      "00011111101000000000000000000011", --  179 -  716
      "00100000000111010000000000111100", --  180 -  720
      "00010000000000000000000000000010", --  181 -  724
      "00100000000111010000000000000000", --  182 -  728
      "00010100101100110000000001001010", --  183 -  732
      "10101111101001010000010101000100", --  184 -  736
      "10001100000111010000010110101100", --  185 -  740
      "00011111101000000000000000000011", --  186 -  744
      "00100000000111010000000000111100", --  187 -  748
      "00010000000000000000000000000010", --  188 -  752
      "00100000000111010000000000000000", --  189 -  756
      "00010100110101000000000001000011", --  190 -  760
      "10101111101001100000010101001000", --  191 -  764
      "10001100000111010000010110101100", --  192 -  768
      "00011111101000000000000000000011", --  193 -  772
      "00100000000111010000000000111100", --  194 -  776
      "00010000000000000000000000000010", --  195 -  780
      "00100000000111010000000000000000", --  196 -  784
      "00010100111101010000000000111100", --  197 -  788
      "10101111101001110000010101001100", --  198 -  792
      "10001100000111010000010110101100", --  199 -  796
      "00011111101000000000000000000011", --  200 -  800
      "00100000000111010000000000111100", --  201 -  804
      "00010000000000000000000000000010", --  202 -  808
      "00100000000111010000000000000000", --  203 -  812
      "00010101000101100000000000110101", --  204 -  816
      "10101111101010000000010101010000", --  205 -  820
      "10001100000111010000010110101100", --  206 -  824
      "00011111101000000000000000000011", --  207 -  828
      "00100000000111010000000000111100", --  208 -  832
      "00010000000000000000000000000010", --  209 -  836
      "00100000000111010000000000000000", --  210 -  840
      "00010101001101110000000000101110", --  211 -  844
      "10101111101010010000010101010100", --  212 -  848
      "10001100000111010000010110101100", --  213 -  852
      "00011111101000000000000000000011", --  214 -  856
      "00100000000111010000000000111100", --  215 -  860
      "00010000000000000000000000000010", --  216 -  864
      "00100000000111010000000000000000", --  217 -  868
      "00010101010110000000000000100111", --  218 -  872
      "10101111101010100000010101011000", --  219 -  876
      "10001100000111010000010110101100", --  220 -  880
      "00011111101000000000000000000011", --  221 -  884
      "00100000000111010000000000111100", --  222 -  888
      "00010000000000000000000000000010", --  223 -  892
      "00100000000111010000000000000000", --  224 -  896
      "00010101011110010000000000100000", --  225 -  900
      "10101111101010110000010101011100", --  226 -  904
      "10001100000111010000010110101100", --  227 -  908
      "00011111101000000000000000000011", --  228 -  912
      "00100000000111010000000000111100", --  229 -  916
      "00010000000000000000000000000010", --  230 -  920
      "00100000000111010000000000000000", --  231 -  924
      "00010101100110100000000000011001", --  232 -  928
      "10101111101011000000010101100000", --  233 -  932
      "10001100000111010000010110101100", --  234 -  936
      "00011111101000000000000000000011", --  235 -  940
      "00100000000111010000000000111100", --  236 -  944
      "00010000000000000000000000000010", --  237 -  948
      "00100000000111010000000000000000", --  238 -  952
      "00010101101110110000000000010010", --  239 -  956
      "10101111101011010000010101100100", --  240 -  960
      "10001100000111010000010110101100", --  241 -  964
      "00011111101000000000000000000011", --  242 -  968
      "00100000000111010000000000111100", --  243 -  972
      "00010000000000000000000000000010", --  244 -  976
      "00100000000111010000000000000000", --  245 -  980
      "00010101110111000000000000001011", --  246 -  984
      "10101111101011100000010101101000", --  247 -  988
      "10001100000111010000010110101100", --  248 -  992
      "00011111101000000000000000000011", --  249 -  996
      "00100000000111010000000000111100", --  250 - 1000
      "00010000000000000000000000000010", --  251 - 1004
      "00100000000111010000000000000000", --  252 - 1008
      "00010111110111110000000000000100", --  253 - 1012
      "10101111101111100000010101101100", --  254 - 1016
      "10101100000111010000010110101100", --  255 - 1020
      "00010000000000001111111110001010", --  256 - 1024
      "10001100000111010000010110101100", --  257 - 1028
      "10001111101000010000010100110100", --  258 - 1032
      "10001100000111010000010110101100", --  259 - 1036
      "10001111101011110000010100110100", --  260 - 1040
      "00010100001011111111111111111100", --  261 - 1044
      "10001100000111010000010110101100", --  262 - 1048
      "10001111101000100000010100111000", --  263 - 1052
      "10001100000111010000010110101100", --  264 - 1056
      "10001111101100000000010100111000", --  265 - 1060
      "00010100010100001111111111111100", --  266 - 1064
      "10001100000111010000010110101100", --  267 - 1068
      "10001111101000110000010100111100", --  268 - 1072
      "10001100000111010000010110101100", --  269 - 1076
      "10001111101100010000010100111100", --  270 - 1080
      "00010100011100011111111111111100", --  271 - 1084
      "10001100000111010000010110101100", --  272 - 1088
      "10001111101001000000010101000000", --  273 - 1092
      "10001100000111010000010110101100", --  274 - 1096
      "10001111101100100000010101000000", --  275 - 1100
      "00010100100100101111111111111100", --  276 - 1104
      "10001100000111010000010110101100", --  277 - 1108
      "10001111101001010000010101000100", --  278 - 1112
      "10001100000111010000010110101100", --  279 - 1116
      "10001111101100110000010101000100", --  280 - 1120
      "00010100101100111111111111111100", --  281 - 1124
      "10001100000111010000010110101100", --  282 - 1128
      "10001111101001100000010101001000", --  283 - 1132
      "10001100000111010000010110101100", --  284 - 1136
      "10001111101101000000010101001000", --  285 - 1140
      "00010100110101001111111111111100", --  286 - 1144
      "10001100000111010000010110101100", --  287 - 1148
      "10001111101001110000010101001100", --  288 - 1152
      "10001100000111010000010110101100", --  289 - 1156
      "10001111101101010000010101001100", --  290 - 1160
      "00010100111101011111111111111100", --  291 - 1164
      "10001100000111010000010110101100", --  292 - 1168
      "10001111101010000000010101010000", --  293 - 1172
      "10001100000111010000010110101100", --  294 - 1176
      "10001111101101100000010101010000", --  295 - 1180
      "00010101000101101111111111111100", --  296 - 1184
      "10001100000111010000010110101100", --  297 - 1188
      "10001111101010010000010101010100", --  298 - 1192
      "10001100000111010000010110101100", --  299 - 1196
      "10001111101101110000010101010100", --  300 - 1200
      "00010101001101111111111111111100", --  301 - 1204
      "10001100000111010000010110101100", --  302 - 1208
      "10001111101010100000010101011000", --  303 - 1212
      "10001100000111010000010110101100", --  304 - 1216
      "10001111101110000000010101011000", --  305 - 1220
      "00010101010110001111111111111100", --  306 - 1224
      "10001100000111010000010110101100", --  307 - 1228
      "10001111101010110000010101011100", --  308 - 1232
      "10001100000111010000010110101100", --  309 - 1236
      "10001111101110010000010101011100", --  310 - 1240
      "00010101011110011111111111111100", --  311 - 1244
      "10001100000111010000010110101100", --  312 - 1248
      "10001111101011000000010101100000", --  313 - 1252
      "10001100000111010000010110101100", --  314 - 1256
      "10001111101110100000010101100000", --  315 - 1260
      "00010101100110101111111111111100", --  316 - 1264
      "10001100000111010000010110101100", --  317 - 1268
      "10001111101011010000010101100100", --  318 - 1272
      "10001100000111010000010110101100", --  319 - 1276
      "10001111101110110000010101100100", --  320 - 1280
      "00010101101110111111111111111100", --  321 - 1284
      "10001100000111010000010110101100", --  322 - 1288
      "10001111101011100000010101101000", --  323 - 1292
      "10001100000111010000010110101100", --  324 - 1296
      "10001111101111000000010101101000", --  325 - 1300
      "00010101110111001111111111111100", --  326 - 1304
      "10001100000111010000010110101100", --  327 - 1308
      "10001111101111100000010101101100", --  328 - 1312
      "10001100000111010000010110101100", --  329 - 1316
      "10001111101111110000010101101100", --  330 - 1320
      "00010111110111111111111111111100", --  331 - 1324
      "00010000000000001111111100111110", --  332 - 1328
      "00000000000000000000000000000000", --  333 - 1332
      "00000000000000000000000000000000", --  334 - 1336
      "00000000000000000000000000000000", --  335 - 1340
      "00000000000000000000000000000000", --  336 - 1344
      "00000000000000000000000000000000", --  337 - 1348
      "00000000000000000000000000000000", --  338 - 1352
      "00000000000000000000000000000000", --  339 - 1356
      "00000000000000000000000000000000", --  340 - 1360
      "00000000000000000000000000000000", --  341 - 1364
      "00000000000000000000000000000000", --  342 - 1368
      "00000000000000000000000000000000", --  343 - 1372
      "00000000000000000000000000000000", --  344 - 1376
      "00000000000000000000000000000000", --  345 - 1380
      "00000000000000000000000000000000", --  346 - 1384
      "00000000000000000000000000000000", --  347 - 1388
      "00000000000000000000000000000000", --  348 - 1392
      "00000000000000000000000000000000", --  349 - 1396
      "00000000000000000000000000000000", --  350 - 1400
      "00000000000000000000000000000000", --  351 - 1404
      "00000000000000000000000000000000", --  352 - 1408
      "00000000000000000000000000000000", --  353 - 1412
      "00000000000000000000000000000000", --  354 - 1416
      "00000000000000000000000000000000", --  355 - 1420
      "00000000000000000000000000000000", --  356 - 1424
      "00000000000000000000000000000000", --  357 - 1428
      "00000000000000000000000000000000", --  358 - 1432
      "00000000000000000000000000000000", --  359 - 1436
      "00000000000000000000000000000000", --  360 - 1440
      "00000000000000000000000000000000", --  361 - 1444
      "00000000000000000000000000000000", --  362 - 1448
      "00000000000000000000001111100111", --  363 - 1452
      "00000000000000000000000000000000", --  364 - 1456
      "00000000000000000000000000000000", --  365 - 1460
      "00000000000000000000000000000000", --  366 - 1464
      "00000000000000000000000000000000", --  367 - 1468
      "00000000000000000000000000000000", --  368 - 1472
      "00000000000000000000000000000000", --  369 - 1476
      "00000000000000000000000000000000", --  370 - 1480
      "00000000000000000000000000000000", --  371 - 1484
      "00000000000000000000000000000000", --  372 - 1488
      "00000000000000000000000000000000", --  373 - 1492
      "00000000000000000000000000000000", --  374 - 1496
      "00000000000000000000000000000000", --  375 - 1500
      "00000000000000000000000000000000", --  376 - 1504
      "00000000000000000000000000000000", --  377 - 1508
      "00000000000000000000000000000000", --  378 - 1512
      "00000000000000000000000000000000", --  379 - 1516
      "00000000000000000000000000000000", --  380 - 1520
      "00000000000000000000000000000000", --  381 - 1524
      "00000000000000000000000000000000", --  382 - 1528
      "00000000000000000000000000000000", --  383 - 1532
      "00000000000000000000000000000000", --  384 - 1536
      "00000000000000000000000000000000", --  385 - 1540
      "00000000000000000000000000000000", --  386 - 1544
      "00000000000000000000000000000000", --  387 - 1548
      "00000000000000000000000000000000", --  388 - 1552
      "00000000000000000000000000000000", --  389 - 1556
      "00000000000000000000000000000000", --  390 - 1560
      "00000000000000000000000000000000", --  391 - 1564
      "00000000000000000000000000000000", --  392 - 1568
      "00000000000000000000000000000000", --  393 - 1572
      "00000000000000000000000000000000", --  394 - 1576
      "00000000000000000000000000000000", --  395 - 1580
      "00000000000000000000000000000000", --  396 - 1584
      "00000000000000000000000000000000", --  397 - 1588
      "00000000000000000000000000000000");--  398 - 1592

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000011101010000101101";
         f_reg(4) <= "00000000000000000001010011000011";
         f_reg(5) <= "00000000000000100001110111000000";
         f_reg(6) <= "00111000001001000010001100100111";
         f_reg(7) <= "00000000001001000010100000100101";
         f_reg(8) <= "00111000010001100000110100110100";
         f_reg(9) <= "00101100011001110100011001001000";
         f_reg(10) <= "00100100110010001111010001101010";
         f_reg(11) <= "00000000110001010100100000000110";
         f_reg(12) <= "00100001000010101000111000000001";
         f_reg(13) <= "00000000000001010101100000000111";
         f_reg(14) <= "00000000110001100110000000000100";
         f_reg(15) <= "00110101001011010100110100111001";
         f_reg(16) <= "00000000000011000111000010000011";
         f_reg(17) <= "10101100000000100000001000111100";
         f_reg(18) <= "00110001110011110111100111000111";
         f_reg(19) <= "00000000000000000000000000000000";
         f_reg(20) <= "00000000000000000000000000000000";
         f_reg(21) <= "00101001001100001101011001101000";
         f_reg(22) <= "10101100000001110000001001000000";
         f_reg(23) <= "00000000000010111000110111000010";
         f_reg(24) <= "00100110001100101011010101001001";
         f_reg(25) <= "00000000000000000000000000000000";
         f_reg(26) <= "00111100000100111000101011001111";
         f_reg(27) <= "00000000000000000000000000000000";
         f_reg(28) <= "00000000000100111010010101000010";
         f_reg(29) <= "00000001101101001010100000100011";
         f_reg(30) <= "00110100011101100011000000000110";
         f_reg(31) <= "10101100000010100000001001000100";
         f_reg(32) <= "00100110000101111111011111011000";
         f_reg(33) <= "00000000000101111100000110000011";
         f_reg(34) <= "00000000000000000000000000000000";
         f_reg(35) <= "10101100000101100000001001001000";
         f_reg(36) <= "00000010101110001100100000100111";
         f_reg(37) <= "00000000000000000000000000000000";
         f_reg(38) <= "10101100000011110000001001001100";
         f_reg(39) <= "00000010010110011101000000101011";
         f_reg(40) <= "00000000000000000000000000000000";
         f_reg(41) <= "10101100000100010000001001010000";
         f_reg(42) <= "00000000000000000000000000000000";
         f_reg(43) <= "10101100000110100000001001010100";
         f_reg(44) <= "00100011111111111111111111111111";
         f_reg(45) <= "00011111111000001111111111010110";
         f_reg(46) <= "00010000000000000000000101100001";
         f_reg(47) <= "00111100000111100000001111100111";
         f_reg(48) <= "00111100000111110000001111100111";
         f_reg(49) <= "00000000000111101111010000000010";
         f_reg(50) <= "00000000000111111111110000000010";
         f_reg(51) <= "00111100000000011101010000101101";
         f_reg(52) <= "00111100000011111101010000101101";
         f_reg(53) <= "00000000000000000001010011000011";
         f_reg(54) <= "00000000000000001000010011000011";
         f_reg(55) <= "00000000000000100001110111000000";
         f_reg(56) <= "00000000000100001000110111000000";
         f_reg(57) <= "00111000001001000010001100100111";
         f_reg(58) <= "00111001111100100010001100100111";
         f_reg(59) <= "00000000001001000010100000100101";
         f_reg(60) <= "00000001111100101001100000100101";
         f_reg(61) <= "00111000010001100000110100110100";
         f_reg(62) <= "00111010000101000000110100110100";
         f_reg(63) <= "00101100011001110100011001001000";
         f_reg(64) <= "00101110001101010100011001001000";
         f_reg(65) <= "00100100110010001111010001101010";
         f_reg(66) <= "00100110100101101111010001101010";
         f_reg(67) <= "00000000110001010100100000000110";
         f_reg(68) <= "00000010100100111011100000000110";
         f_reg(69) <= "00100001000010101000111000000001";
         f_reg(70) <= "00100010110110001000111000000001";
         f_reg(71) <= "00000000000001010101100000000111";
         f_reg(72) <= "00000000000100111100100000000111";
         f_reg(73) <= "00000000110001100110000000000100";
         f_reg(74) <= "00000010100101001101000000000100";
         f_reg(75) <= "00110101001011010100110100111001";
         f_reg(76) <= "00110110111110110100110100111001";
         f_reg(77) <= "00000000000011000111000010000011";
         f_reg(78) <= "00000000000110101110000010000011";
         f_reg(79) <= "00010100010100000000000010110011";
         f_reg(80) <= "10101100000000100000001000111100";
         f_reg(81) <= "00110001110000010111100111000111";
         f_reg(82) <= "00110011100011110111100111000111";
         f_reg(83) <= "00000000000000000000000000000000";
         f_reg(84) <= "00000000000000000000000000000000";
         f_reg(85) <= "00000000000000000000000000000000";
         f_reg(86) <= "00000000000000000000000000000000";
         f_reg(87) <= "00101001001001001101011001101000";
         f_reg(88) <= "00101010111100101101011001101000";
         f_reg(89) <= "00010100111101010000000010101001";
         f_reg(90) <= "10101100000001110000001001000000";
         f_reg(91) <= "00000000000010110100010111000010";
         f_reg(92) <= "00000000000110011011010111000010";
         f_reg(93) <= "00100101000001011011010101001001";
         f_reg(94) <= "00100110110100111011010101001001";
         f_reg(95) <= "00000000000000000000000000000000";
         f_reg(96) <= "00000000000000000000000000000000";
         f_reg(97) <= "00111100000001101000101011001111";
         f_reg(98) <= "00111100000101001000101011001111";
         f_reg(99) <= "00000000000000000000000000000000";
         f_reg(100) <= "00000000000000000000000000000000";
         f_reg(101) <= "00000000000001100110010101000010";
         f_reg(102) <= "00000000000101001101010101000010";
         f_reg(103) <= "00000001101011000001000000100011";
         f_reg(104) <= "00000011011110101000000000100011";
         f_reg(105) <= "00110100011011100011000000000110";
         f_reg(106) <= "00110110001111000011000000000110";
         f_reg(107) <= "00010101010110000000000010010111";
         f_reg(108) <= "10101100000010100000001001000100";
         f_reg(109) <= "00100100100010011111011111011000";
         f_reg(110) <= "00100110010101111111011111011000";
         f_reg(111) <= "00000000000010010011100110000011";
         f_reg(112) <= "00000000000101111010100110000011";
         f_reg(113) <= "00000000000000000000000000000000";
         f_reg(114) <= "00000000000000000000000000000000";
         f_reg(115) <= "00010101110111000000000010001111";
         f_reg(116) <= "10101100000011100000001001001000";
         f_reg(117) <= "00000000010001110101100000100111";
         f_reg(118) <= "00000010000101011100100000100111";
         f_reg(119) <= "00000000000000000000000000000000";
         f_reg(120) <= "00000000000000000000000000000000";
         f_reg(121) <= "00010100001011110000000010001001";
         f_reg(122) <= "10101100000000010000001001001100";
         f_reg(123) <= "00000000101010110011000000101011";
         f_reg(124) <= "00000010011110011010000000101011";
         f_reg(125) <= "00000000000000000000000000000000";
         f_reg(126) <= "00000000000000000000000000000000";
         f_reg(127) <= "00010101000101100000000010000011";
         f_reg(128) <= "10101100000010000000001001010000";
         f_reg(129) <= "00000000000000000000000000000000";
         f_reg(130) <= "00000000000000000000000000000000";
         f_reg(131) <= "00010100110101000000000001111111";
         f_reg(132) <= "10101100000001100000001001010100";
         f_reg(133) <= "00100011110111011111111100000110";
         f_reg(134) <= "00010011101000000000000000010001";
         f_reg(135) <= "00100011110111011111111000001100";
         f_reg(136) <= "00010011101000000000000000001111";
         f_reg(137) <= "00100011110111011111110100010010";
         f_reg(138) <= "00010011101000000000000000001101";
         f_reg(139) <= "00100011110111101111111111111111";
         f_reg(140) <= "00100011111111111111111111111111";
         f_reg(141) <= "00010111110111110000000001110101";
         f_reg(142) <= "00011111111000001111111110100101";
         f_reg(143) <= "00010000000000000000000100000000";
         f_reg(144) <= "00000000000000000000000000000000";
         f_reg(145) <= "00000000000000000000000000000000";
         f_reg(146) <= "00000000000000000000000000000000";
         f_reg(147) <= "00000000000000000000000000000000";
         f_reg(148) <= "00000000000000000000000000000000";
         f_reg(149) <= "00000000000000000000000000000000";
         f_reg(150) <= "00000000000000000000000000000000";
         f_reg(151) <= "10001100000111010000010110101100";
         f_reg(152) <= "00011111101000000000000000000011";
         f_reg(153) <= "00100000000111010000000000111100";
         f_reg(154) <= "00010000000000000000000000000010";
         f_reg(155) <= "00100000000111010000000000000000";
         f_reg(156) <= "00010100001011110000000001100110";
         f_reg(157) <= "10101111101000010000010100110100";
         f_reg(158) <= "10001100000111010000010110101100";
         f_reg(159) <= "00011111101000000000000000000011";
         f_reg(160) <= "00100000000111010000000000111100";
         f_reg(161) <= "00010000000000000000000000000010";
         f_reg(162) <= "00100000000111010000000000000000";
         f_reg(163) <= "00010100010100000000000001011111";
         f_reg(164) <= "10101111101000100000010100111000";
         f_reg(165) <= "10001100000111010000010110101100";
         f_reg(166) <= "00011111101000000000000000000011";
         f_reg(167) <= "00100000000111010000000000111100";
         f_reg(168) <= "00010000000000000000000000000010";
         f_reg(169) <= "00100000000111010000000000000000";
         f_reg(170) <= "00010100011100010000000001011000";
         f_reg(171) <= "10101111101000110000010100111100";
         f_reg(172) <= "10001100000111010000010110101100";
         f_reg(173) <= "00011111101000000000000000000011";
         f_reg(174) <= "00100000000111010000000000111100";
         f_reg(175) <= "00010000000000000000000000000010";
         f_reg(176) <= "00100000000111010000000000000000";
         f_reg(177) <= "00010100100100100000000001010001";
         f_reg(178) <= "10101111101001000000010101000000";
         f_reg(179) <= "10001100000111010000010110101100";
         f_reg(180) <= "00011111101000000000000000000011";
         f_reg(181) <= "00100000000111010000000000111100";
         f_reg(182) <= "00010000000000000000000000000010";
         f_reg(183) <= "00100000000111010000000000000000";
         f_reg(184) <= "00010100101100110000000001001010";
         f_reg(185) <= "10101111101001010000010101000100";
         f_reg(186) <= "10001100000111010000010110101100";
         f_reg(187) <= "00011111101000000000000000000011";
         f_reg(188) <= "00100000000111010000000000111100";
         f_reg(189) <= "00010000000000000000000000000010";
         f_reg(190) <= "00100000000111010000000000000000";
         f_reg(191) <= "00010100110101000000000001000011";
         f_reg(192) <= "10101111101001100000010101001000";
         f_reg(193) <= "10001100000111010000010110101100";
         f_reg(194) <= "00011111101000000000000000000011";
         f_reg(195) <= "00100000000111010000000000111100";
         f_reg(196) <= "00010000000000000000000000000010";
         f_reg(197) <= "00100000000111010000000000000000";
         f_reg(198) <= "00010100111101010000000000111100";
         f_reg(199) <= "10101111101001110000010101001100";
         f_reg(200) <= "10001100000111010000010110101100";
         f_reg(201) <= "00011111101000000000000000000011";
         f_reg(202) <= "00100000000111010000000000111100";
         f_reg(203) <= "00010000000000000000000000000010";
         f_reg(204) <= "00100000000111010000000000000000";
         f_reg(205) <= "00010101000101100000000000110101";
         f_reg(206) <= "10101111101010000000010101010000";
         f_reg(207) <= "10001100000111010000010110101100";
         f_reg(208) <= "00011111101000000000000000000011";
         f_reg(209) <= "00100000000111010000000000111100";
         f_reg(210) <= "00010000000000000000000000000010";
         f_reg(211) <= "00100000000111010000000000000000";
         f_reg(212) <= "00010101001101110000000000101110";
         f_reg(213) <= "10101111101010010000010101010100";
         f_reg(214) <= "10001100000111010000010110101100";
         f_reg(215) <= "00011111101000000000000000000011";
         f_reg(216) <= "00100000000111010000000000111100";
         f_reg(217) <= "00010000000000000000000000000010";
         f_reg(218) <= "00100000000111010000000000000000";
         f_reg(219) <= "00010101010110000000000000100111";
         f_reg(220) <= "10101111101010100000010101011000";
         f_reg(221) <= "10001100000111010000010110101100";
         f_reg(222) <= "00011111101000000000000000000011";
         f_reg(223) <= "00100000000111010000000000111100";
         f_reg(224) <= "00010000000000000000000000000010";
         f_reg(225) <= "00100000000111010000000000000000";
         f_reg(226) <= "00010101011110010000000000100000";
         f_reg(227) <= "10101111101010110000010101011100";
         f_reg(228) <= "10001100000111010000010110101100";
         f_reg(229) <= "00011111101000000000000000000011";
         f_reg(230) <= "00100000000111010000000000111100";
         f_reg(231) <= "00010000000000000000000000000010";
         f_reg(232) <= "00100000000111010000000000000000";
         f_reg(233) <= "00010101100110100000000000011001";
         f_reg(234) <= "10101111101011000000010101100000";
         f_reg(235) <= "10001100000111010000010110101100";
         f_reg(236) <= "00011111101000000000000000000011";
         f_reg(237) <= "00100000000111010000000000111100";
         f_reg(238) <= "00010000000000000000000000000010";
         f_reg(239) <= "00100000000111010000000000000000";
         f_reg(240) <= "00010101101110110000000000010010";
         f_reg(241) <= "10101111101011010000010101100100";
         f_reg(242) <= "10001100000111010000010110101100";
         f_reg(243) <= "00011111101000000000000000000011";
         f_reg(244) <= "00100000000111010000000000111100";
         f_reg(245) <= "00010000000000000000000000000010";
         f_reg(246) <= "00100000000111010000000000000000";
         f_reg(247) <= "00010101110111000000000000001011";
         f_reg(248) <= "10101111101011100000010101101000";
         f_reg(249) <= "10001100000111010000010110101100";
         f_reg(250) <= "00011111101000000000000000000011";
         f_reg(251) <= "00100000000111010000000000111100";
         f_reg(252) <= "00010000000000000000000000000010";
         f_reg(253) <= "00100000000111010000000000000000";
         f_reg(254) <= "00010111110111110000000000000100";
         f_reg(255) <= "10101111101111100000010101101100";
         f_reg(256) <= "10101100000111010000010110101100";
         f_reg(257) <= "00010000000000001111111110001010";
         f_reg(258) <= "10001100000111010000010110101100";
         f_reg(259) <= "10001111101000010000010100110100";
         f_reg(260) <= "10001100000111010000010110101100";
         f_reg(261) <= "10001111101011110000010100110100";
         f_reg(262) <= "00010100001011111111111111111100";
         f_reg(263) <= "10001100000111010000010110101100";
         f_reg(264) <= "10001111101000100000010100111000";
         f_reg(265) <= "10001100000111010000010110101100";
         f_reg(266) <= "10001111101100000000010100111000";
         f_reg(267) <= "00010100010100001111111111111100";
         f_reg(268) <= "10001100000111010000010110101100";
         f_reg(269) <= "10001111101000110000010100111100";
         f_reg(270) <= "10001100000111010000010110101100";
         f_reg(271) <= "10001111101100010000010100111100";
         f_reg(272) <= "00010100011100011111111111111100";
         f_reg(273) <= "10001100000111010000010110101100";
         f_reg(274) <= "10001111101001000000010101000000";
         f_reg(275) <= "10001100000111010000010110101100";
         f_reg(276) <= "10001111101100100000010101000000";
         f_reg(277) <= "00010100100100101111111111111100";
         f_reg(278) <= "10001100000111010000010110101100";
         f_reg(279) <= "10001111101001010000010101000100";
         f_reg(280) <= "10001100000111010000010110101100";
         f_reg(281) <= "10001111101100110000010101000100";
         f_reg(282) <= "00010100101100111111111111111100";
         f_reg(283) <= "10001100000111010000010110101100";
         f_reg(284) <= "10001111101001100000010101001000";
         f_reg(285) <= "10001100000111010000010110101100";
         f_reg(286) <= "10001111101101000000010101001000";
         f_reg(287) <= "00010100110101001111111111111100";
         f_reg(288) <= "10001100000111010000010110101100";
         f_reg(289) <= "10001111101001110000010101001100";
         f_reg(290) <= "10001100000111010000010110101100";
         f_reg(291) <= "10001111101101010000010101001100";
         f_reg(292) <= "00010100111101011111111111111100";
         f_reg(293) <= "10001100000111010000010110101100";
         f_reg(294) <= "10001111101010000000010101010000";
         f_reg(295) <= "10001100000111010000010110101100";
         f_reg(296) <= "10001111101101100000010101010000";
         f_reg(297) <= "00010101000101101111111111111100";
         f_reg(298) <= "10001100000111010000010110101100";
         f_reg(299) <= "10001111101010010000010101010100";
         f_reg(300) <= "10001100000111010000010110101100";
         f_reg(301) <= "10001111101101110000010101010100";
         f_reg(302) <= "00010101001101111111111111111100";
         f_reg(303) <= "10001100000111010000010110101100";
         f_reg(304) <= "10001111101010100000010101011000";
         f_reg(305) <= "10001100000111010000010110101100";
         f_reg(306) <= "10001111101110000000010101011000";
         f_reg(307) <= "00010101010110001111111111111100";
         f_reg(308) <= "10001100000111010000010110101100";
         f_reg(309) <= "10001111101010110000010101011100";
         f_reg(310) <= "10001100000111010000010110101100";
         f_reg(311) <= "10001111101110010000010101011100";
         f_reg(312) <= "00010101011110011111111111111100";
         f_reg(313) <= "10001100000111010000010110101100";
         f_reg(314) <= "10001111101011000000010101100000";
         f_reg(315) <= "10001100000111010000010110101100";
         f_reg(316) <= "10001111101110100000010101100000";
         f_reg(317) <= "00010101100110101111111111111100";
         f_reg(318) <= "10001100000111010000010110101100";
         f_reg(319) <= "10001111101011010000010101100100";
         f_reg(320) <= "10001100000111010000010110101100";
         f_reg(321) <= "10001111101110110000010101100100";
         f_reg(322) <= "00010101101110111111111111111100";
         f_reg(323) <= "10001100000111010000010110101100";
         f_reg(324) <= "10001111101011100000010101101000";
         f_reg(325) <= "10001100000111010000010110101100";
         f_reg(326) <= "10001111101111000000010101101000";
         f_reg(327) <= "00010101110111001111111111111100";
         f_reg(328) <= "10001100000111010000010110101100";
         f_reg(329) <= "10001111101111100000010101101100";
         f_reg(330) <= "10001100000111010000010110101100";
         f_reg(331) <= "10001111101111110000010101101100";
         f_reg(332) <= "00010111110111111111111111111100";
         f_reg(333) <= "00010000000000001111111100111110";
         f_reg(334) <= "00000000000000000000000000000000";
         f_reg(335) <= "00000000000000000000000000000000";
         f_reg(336) <= "00000000000000000000000000000000";
         f_reg(337) <= "00000000000000000000000000000000";
         f_reg(338) <= "00000000000000000000000000000000";
         f_reg(339) <= "00000000000000000000000000000000";
         f_reg(340) <= "00000000000000000000000000000000";
         f_reg(341) <= "00000000000000000000000000000000";
         f_reg(342) <= "00000000000000000000000000000000";
         f_reg(343) <= "00000000000000000000000000000000";
         f_reg(344) <= "00000000000000000000000000000000";
         f_reg(345) <= "00000000000000000000000000000000";
         f_reg(346) <= "00000000000000000000000000000000";
         f_reg(347) <= "00000000000000000000000000000000";
         f_reg(348) <= "00000000000000000000000000000000";
         f_reg(349) <= "00000000000000000000000000000000";
         f_reg(350) <= "00000000000000000000000000000000";
         f_reg(351) <= "00000000000000000000000000000000";
         f_reg(352) <= "00000000000000000000000000000000";
         f_reg(353) <= "00000000000000000000000000000000";
         f_reg(354) <= "00000000000000000000000000000000";
         f_reg(355) <= "00000000000000000000000000000000";
         f_reg(356) <= "00000000000000000000000000000000";
         f_reg(357) <= "00000000000000000000000000000000";
         f_reg(358) <= "00000000000000000000000000000000";
         f_reg(359) <= "00000000000000000000000000000000";
         f_reg(360) <= "00000000000000000000000000000000";
         f_reg(361) <= "00000000000000000000000000000000";
         f_reg(362) <= "00000000000000000000000000000000";
         f_reg(363) <= "00000000000000000000000000000000";
         f_reg(364) <= "00000000000000000000001111100111";
         f_reg(365) <= "00000000000000000000000000000000";
         f_reg(366) <= "00000000000000000000000000000000";
         f_reg(367) <= "00000000000000000000000000000000";
         f_reg(368) <= "00000000000000000000000000000000";
         f_reg(369) <= "00000000000000000000000000000000";
         f_reg(370) <= "00000000000000000000000000000000";
         f_reg(371) <= "00000000000000000000000000000000";
         f_reg(372) <= "00000000000000000000000000000000";
         f_reg(373) <= "00000000000000000000000000000000";
         f_reg(374) <= "00000000000000000000000000000000";
         f_reg(375) <= "00000000000000000000000000000000";
         f_reg(376) <= "00000000000000000000000000000000";
         f_reg(377) <= "00000000000000000000000000000000";
         f_reg(378) <= "00000000000000000000000000000000";
         f_reg(379) <= "00000000000000000000000000000000";
         f_reg(380) <= "00000000000000000000000000000000";
         f_reg(381) <= "00000000000000000000000000000000";
         f_reg(382) <= "00000000000000000000000000000000";
         f_reg(383) <= "00000000000000000000000000000000";
         f_reg(384) <= "00000000000000000000000000000000";
         f_reg(385) <= "00000000000000000000000000000000";
         f_reg(386) <= "00000000000000000000000000000000";
         f_reg(387) <= "00000000000000000000000000000000";
         f_reg(388) <= "00000000000000000000000000000000";
         f_reg(389) <= "00000000000000000000000000000000";
         f_reg(390) <= "00000000000000000000000000000000";
         f_reg(391) <= "00000000000000000000000000000000";
         f_reg(392) <= "00000000000000000000000000000000";
         f_reg(393) <= "00000000000000000000000000000000";
         f_reg(394) <= "00000000000000000000000000000000";
         f_reg(395) <= "00000000000000000000000000000000";
         f_reg(396) <= "00000000000000000000000000000000";
         f_reg(397) <= "00000000000000000000000000000000";
         f_reg(398) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 -11219
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SRA R2 R0 19
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SLL R3 R2 23
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- XORI R4 R1 8999
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- OR R5 R1 R4
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- XORI R6 R2 3380
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- SLTIU R7 R3 17992
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- ADDIU R8 R6 -2966
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- SRLV R9 R5 R6
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- ADDI R10 R8 -29183
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- SRAV R11 R5 R0
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- SLLV R12 R6 R6
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- ORI R13 R9 19769
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- SRA R14 R12 2
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- SW R2 R0 572
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- ANDI R15 R14 31175
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- NOP
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- NOP
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SLTI R16 R9 -10648
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- SW R7 R0 576
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- SRL R17 R11 23
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- ADDIU R18 R17 -19127
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- NOP
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- LUI R19 -30001
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- NOP
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- SRL R20 R19 21
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- SUBU R21 R13 R20
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- ORI R22 R3 12294
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- SW R10 R0 580
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- ADDIU R23 R16 -2088
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- SRA R24 R23 6
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- NOP
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- SW R22 R0 584
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- NOR R25 R21 R24
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- NOP
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- SW R15 R0 588
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- SLTU R26 R18 R25
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- NOP
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- SW R17 R0 592
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- NOP
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SW R26 R0 596
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- BGTZ R31 -42
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- BEQ R0 R0 353
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- LUI R30 999
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- LUI R31 999
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- LUI R1 -11219
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- LUI R15 -11219
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- SRA R2 R0 19
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SRA R16 R0 19
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SLL R3 R2 23
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- SLL R17 R16 23
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- XORI R4 R1 8999
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- XORI R18 R15 8999
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- OR R5 R1 R4
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- OR R19 R15 R18
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- XORI R6 R2 3380
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- XORI R20 R16 3380
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- SLTIU R7 R3 17992
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- SLTIU R21 R17 17992
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- ADDIU R8 R6 -2966
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- ADDIU R22 R20 -2966
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- SRLV R9 R5 R6
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- SRLV R23 R19 R20
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- ADDI R10 R8 -29183
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- ADDI R24 R22 -29183
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- SRAV R11 R5 R0
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- SRAV R25 R19 R0
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SLLV R12 R6 R6
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- SLLV R26 R20 R20
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- ORI R13 R9 19769
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- ORI R27 R23 19769
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- SRA R14 R12 2
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- SRA R28 R26 2
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- BNE R2 R16 179
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- SW R2 R0 572
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- ANDI R1 R14 31175
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- ANDI R15 R28 31175
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- NOP
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- NOP
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- NOP
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- NOP
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SLTI R4 R9 -10648
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- SLTI R18 R23 -10648
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- BNE R7 R21 169
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- SW R7 R0 576
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- SRL R8 R11 23
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- SRL R22 R25 23
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- ADDIU R5 R8 -19127
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- ADDIU R19 R22 -19127
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- NOP
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- NOP
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- LUI R6 -30001
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- LUI R20 -30001
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- NOP
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- NOP
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- SRL R12 R6 21
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- SRL R26 R20 21
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SUBU R2 R13 R12
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- SUBU R16 R27 R26
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- ORI R14 R3 12294
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- ORI R28 R17 12294
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- BNE R10 R24 151
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- SW R10 R0 580
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- ADDIU R9 R4 -2088
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- ADDIU R23 R18 -2088
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- SRA R7 R9 6
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- SRA R21 R23 6
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- NOP
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- NOP
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- BNE R14 R28 143
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- SW R14 R0 584
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- NOR R11 R2 R7
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- NOR R25 R16 R21
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- NOP
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- NOP
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- BNE R1 R15 137
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- SW R1 R0 588
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- SLTU R6 R5 R11
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SLTU R20 R19 R25
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- NOP
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- NOP
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- BNE R8 R22 131
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SW R8 R0 592
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- NOP
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- NOP
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- BNE R6 R20 127
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- SW R6 R0 596
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- BEQ R29 R0 17
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- BEQ R29 R0 15
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- BEQ R29 R0 13
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- BNE R30 R31 117
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- BGTZ R31 -91
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- BEQ R0 R0 256
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- NOP
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- NOP
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- NOP
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- NOP
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- NOP
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- NOP
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- NOP
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- SW R1 R29 1332
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- SW R2 R29 1336
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- SW R3 R29 1340
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- SW R4 R29 1344
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- SW R5 R29 1348
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- SW R6 R29 1352
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- SW R7 R29 1356
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- SW R8 R29 1360
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- SW R9 R29 1364
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- SW R10 R29 1368
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- SW R11 R29 1372
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- SW R12 R29 1376
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- SW R13 R29 1380
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- SW R14 R29 1384
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- SW R30 R29 1388
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- SW R29 R0 1452
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- BEQ R0 R0 -118
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- LW R1 R29 1332
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- LW R15 R29 1332
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- LW R2 R29 1336
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- LW R16 R29 1336
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- LW R3 R29 1340
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- LW R17 R29 1340
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- LW R4 R29 1344
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- LW R18 R29 1344
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- LW R5 R29 1348
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- LW R19 R29 1348
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- LW R6 R29 1352
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- LW R20 R29 1352
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- LW R7 R29 1356
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- LW R21 R29 1356
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- LW R8 R29 1360
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- LW R22 R29 1360
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- LW R9 R29 1364
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- LW R23 R29 1364
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- LW R10 R29 1368
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- LW R24 R29 1368
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- LW R11 R29 1372
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- LW R25 R29 1372
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- LW R12 R29 1376
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- LW R26 R29 1376
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- LW R13 R29 1380
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- LW R27 R29 1380
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- LW R14 R29 1384
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- LW R28 R29 1384
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- LW R30 R29 1388
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- LW R29 R0 1452
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- LW R31 R29 1388
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- BEQ R0 R0 -194
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- NOP
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- NOP
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- NOP
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- NOP
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- NOP
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- NOP
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- NOP
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- NOP
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- NOP
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- NOP
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- NOP
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- NOP
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- NOP
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- NOP
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- NOP
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- NOP
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- NOP
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- NOP
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- NOP
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- NOP
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- NOP
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- NOP
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- NOP
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- NOP
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- NOP
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- NOP
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- NOP
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- NOP
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- NOP
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- NOP
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- NOP
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- NOP
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- NOP
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- NOP
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- NOP
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- NOP
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- NOP
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- NOP
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- NOP
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- NOP
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- NOP
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- NOP
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- NOP
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- NOP
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- NOP
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- NOP
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- NOP
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- NOP
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- NOP
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- NOP
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- NOP
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- NOP
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- NOP
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- NOP
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- NOP
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- NOP
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- NOP
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- NOP
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- NOP
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- NOP
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- NOP
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- NOP
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- NOP
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- NOP
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- NOP
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011101010000101101";
                        f_reg(4) <= "00000000000000000001010011000011";
                        f_reg(5) <= "00000000000000100001110111000000";
                        f_reg(6) <= "00111000001001000010001100100111";
                        f_reg(7) <= "00000000001001000010100000100101";
                        f_reg(8) <= "00111000010001100000110100110100";
                        f_reg(9) <= "00101100011001110100011001001000";
                        f_reg(10) <= "00100100110010001111010001101010";
                        f_reg(11) <= "00000000110001010100100000000110";
                        f_reg(12) <= "00100001000010101000111000000001";
                        f_reg(13) <= "00000000000001010101100000000111";
                        f_reg(14) <= "00000000110001100110000000000100";
                        f_reg(15) <= "00110101001011010100110100111001";
                        f_reg(16) <= "00000000000011000111000010000011";
                        f_reg(17) <= "10101100000000100000001000111100";
                        f_reg(18) <= "00110001110011110111100111000111";
                        f_reg(19) <= "00000000000000000000000000000000";
                        f_reg(20) <= "00000000000000000000000000000000";
                        f_reg(21) <= "00101001001100001101011001101000";
                        f_reg(22) <= "10101100000001110000001001000000";
                        f_reg(23) <= "00000000000010111000110111000010";
                        f_reg(24) <= "00100110001100101011010101001001";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00111100000100111000101011001111";
                        f_reg(27) <= "00000000000000000000000000000000";
                        f_reg(28) <= "00000000000100111010010101000010";
                        f_reg(29) <= "00000001101101001010100000100011";
                        f_reg(30) <= "00110100011101100011000000000110";
                        f_reg(31) <= "10101100000010100000001001000100";
                        f_reg(32) <= "00100110000101111111011111011000";
                        f_reg(33) <= "00000000000101111100000110000011";
                        f_reg(34) <= "00000000000000000000000000000000";
                        f_reg(35) <= "10101100000101100000001001001000";
                        f_reg(36) <= "00000010101110001100100000100111";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "10101100000011110000001001001100";
                        f_reg(39) <= "00000010010110011101000000101011";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "10101100000100010000001001010000";
                        f_reg(42) <= "00000000000000000000000000000000";
                        f_reg(43) <= "10101100000110100000001001010100";
                        f_reg(44) <= "00100011111111111111111111111111";
                        f_reg(45) <= "00011111111000001111111111010110";
                        f_reg(46) <= "00010000000000000000000101100001";
                        f_reg(47) <= "00111100000111100000001111100111";
                        f_reg(48) <= "00111100000111110000001111100111";
                        f_reg(49) <= "00000000000111101111010000000010";
                        f_reg(50) <= "00000000000111111111110000000010";
                        f_reg(51) <= "00111100000000011101010000101101";
                        f_reg(52) <= "00111100000011111101010000101101";
                        f_reg(53) <= "00000000000000000001010011000011";
                        f_reg(54) <= "00000000000000001000010011000011";
                        f_reg(55) <= "00000000000000100001110111000000";
                        f_reg(56) <= "00000000000100001000110111000000";
                        f_reg(57) <= "00111000001001000010001100100111";
                        f_reg(58) <= "00111001111100100010001100100111";
                        f_reg(59) <= "00000000001001000010100000100101";
                        f_reg(60) <= "00000001111100101001100000100101";
                        f_reg(61) <= "00111000010001100000110100110100";
                        f_reg(62) <= "00111010000101000000110100110100";
                        f_reg(63) <= "00101100011001110100011001001000";
                        f_reg(64) <= "00101110001101010100011001001000";
                        f_reg(65) <= "00100100110010001111010001101010";
                        f_reg(66) <= "00100110100101101111010001101010";
                        f_reg(67) <= "00000000110001010100100000000110";
                        f_reg(68) <= "00000010100100111011100000000110";
                        f_reg(69) <= "00100001000010101000111000000001";
                        f_reg(70) <= "00100010110110001000111000000001";
                        f_reg(71) <= "00000000000001010101100000000111";
                        f_reg(72) <= "00000000000100111100100000000111";
                        f_reg(73) <= "00000000110001100110000000000100";
                        f_reg(74) <= "00000010100101001101000000000100";
                        f_reg(75) <= "00110101001011010100110100111001";
                        f_reg(76) <= "00110110111110110100110100111001";
                        f_reg(77) <= "00000000000011000111000010000011";
                        f_reg(78) <= "00000000000110101110000010000011";
                        f_reg(79) <= "00010100010100000000000010110011";
                        f_reg(80) <= "10101100000000100000001000111100";
                        f_reg(81) <= "00110001110000010111100111000111";
                        f_reg(82) <= "00110011100011110111100111000111";
                        f_reg(83) <= "00000000000000000000000000000000";
                        f_reg(84) <= "00000000000000000000000000000000";
                        f_reg(85) <= "00000000000000000000000000000000";
                        f_reg(86) <= "00000000000000000000000000000000";
                        f_reg(87) <= "00101001001001001101011001101000";
                        f_reg(88) <= "00101010111100101101011001101000";
                        f_reg(89) <= "00010100111101010000000010101001";
                        f_reg(90) <= "10101100000001110000001001000000";
                        f_reg(91) <= "00000000000010110100010111000010";
                        f_reg(92) <= "00000000000110011011010111000010";
                        f_reg(93) <= "00100101000001011011010101001001";
                        f_reg(94) <= "00100110110100111011010101001001";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000000000000000000000000000";
                        f_reg(97) <= "00111100000001101000101011001111";
                        f_reg(98) <= "00111100000101001000101011001111";
                        f_reg(99) <= "00000000000000000000000000000000";
                        f_reg(100) <= "00000000000000000000000000000000";
                        f_reg(101) <= "00000000000001100110010101000010";
                        f_reg(102) <= "00000000000101001101010101000010";
                        f_reg(103) <= "00000001101011000001000000100011";
                        f_reg(104) <= "00000011011110101000000000100011";
                        f_reg(105) <= "00110100011011100011000000000110";
                        f_reg(106) <= "00110110001111000011000000000110";
                        f_reg(107) <= "00010101010110000000000010010111";
                        f_reg(108) <= "10101100000010100000001001000100";
                        f_reg(109) <= "00100100100010011111011111011000";
                        f_reg(110) <= "00100110010101111111011111011000";
                        f_reg(111) <= "00000000000010010011100110000011";
                        f_reg(112) <= "00000000000101111010100110000011";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00010101110111000000000010001111";
                        f_reg(116) <= "10101100000011100000001001001000";
                        f_reg(117) <= "00000000010001110101100000100111";
                        f_reg(118) <= "00000010000101011100100000100111";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000000000000000000000000000";
                        f_reg(121) <= "00010100001011110000000010001001";
                        f_reg(122) <= "10101100000000010000001001001100";
                        f_reg(123) <= "00000000101010110011000000101011";
                        f_reg(124) <= "00000010011110011010000000101011";
                        f_reg(125) <= "00000000000000000000000000000000";
                        f_reg(126) <= "00000000000000000000000000000000";
                        f_reg(127) <= "00010101000101100000000010000011";
                        f_reg(128) <= "10101100000010000000001001010000";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010100110101000000000001111111";
                        f_reg(132) <= "10101100000001100000001001010100";
                        f_reg(133) <= "00100011110111011111111100000110";
                        f_reg(134) <= "00010011101000000000000000010001";
                        f_reg(135) <= "00100011110111011111111000001100";
                        f_reg(136) <= "00010011101000000000000000001111";
                        f_reg(137) <= "00100011110111011111110100010010";
                        f_reg(138) <= "00010011101000000000000000001101";
                        f_reg(139) <= "00100011110111101111111111111111";
                        f_reg(140) <= "00100011111111111111111111111111";
                        f_reg(141) <= "00010111110111110000000001110101";
                        f_reg(142) <= "00011111111000001111111110100101";
                        f_reg(143) <= "00010000000000000000000100000000";
                        f_reg(144) <= "00000000000000000000000000000000";
                        f_reg(145) <= "00000000000000000000000000000000";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000000000000000000000000000";
                        f_reg(149) <= "00000000000000000000000000000000";
                        f_reg(150) <= "00000000000000000000000000000000";
                        f_reg(151) <= "10001100000111010000010110101100";
                        f_reg(152) <= "00011111101000000000000000000011";
                        f_reg(153) <= "00100000000111010000000000111100";
                        f_reg(154) <= "00010000000000000000000000000010";
                        f_reg(155) <= "00100000000111010000000000000000";
                        f_reg(156) <= "00010100001011110000000001100110";
                        f_reg(157) <= "10101111101000010000010100110100";
                        f_reg(158) <= "10001100000111010000010110101100";
                        f_reg(159) <= "00011111101000000000000000000011";
                        f_reg(160) <= "00100000000111010000000000111100";
                        f_reg(161) <= "00010000000000000000000000000010";
                        f_reg(162) <= "00100000000111010000000000000000";
                        f_reg(163) <= "00010100010100000000000001011111";
                        f_reg(164) <= "10101111101000100000010100111000";
                        f_reg(165) <= "10001100000111010000010110101100";
                        f_reg(166) <= "00011111101000000000000000000011";
                        f_reg(167) <= "00100000000111010000000000111100";
                        f_reg(168) <= "00010000000000000000000000000010";
                        f_reg(169) <= "00100000000111010000000000000000";
                        f_reg(170) <= "00010100011100010000000001011000";
                        f_reg(171) <= "10101111101000110000010100111100";
                        f_reg(172) <= "10001100000111010000010110101100";
                        f_reg(173) <= "00011111101000000000000000000011";
                        f_reg(174) <= "00100000000111010000000000111100";
                        f_reg(175) <= "00010000000000000000000000000010";
                        f_reg(176) <= "00100000000111010000000000000000";
                        f_reg(177) <= "00010100100100100000000001010001";
                        f_reg(178) <= "10101111101001000000010101000000";
                        f_reg(179) <= "10001100000111010000010110101100";
                        f_reg(180) <= "00011111101000000000000000000011";
                        f_reg(181) <= "00100000000111010000000000111100";
                        f_reg(182) <= "00010000000000000000000000000010";
                        f_reg(183) <= "00100000000111010000000000000000";
                        f_reg(184) <= "00010100101100110000000001001010";
                        f_reg(185) <= "10101111101001010000010101000100";
                        f_reg(186) <= "10001100000111010000010110101100";
                        f_reg(187) <= "00011111101000000000000000000011";
                        f_reg(188) <= "00100000000111010000000000111100";
                        f_reg(189) <= "00010000000000000000000000000010";
                        f_reg(190) <= "00100000000111010000000000000000";
                        f_reg(191) <= "00010100110101000000000001000011";
                        f_reg(192) <= "10101111101001100000010101001000";
                        f_reg(193) <= "10001100000111010000010110101100";
                        f_reg(194) <= "00011111101000000000000000000011";
                        f_reg(195) <= "00100000000111010000000000111100";
                        f_reg(196) <= "00010000000000000000000000000010";
                        f_reg(197) <= "00100000000111010000000000000000";
                        f_reg(198) <= "00010100111101010000000000111100";
                        f_reg(199) <= "10101111101001110000010101001100";
                        f_reg(200) <= "10001100000111010000010110101100";
                        f_reg(201) <= "00011111101000000000000000000011";
                        f_reg(202) <= "00100000000111010000000000111100";
                        f_reg(203) <= "00010000000000000000000000000010";
                        f_reg(204) <= "00100000000111010000000000000000";
                        f_reg(205) <= "00010101000101100000000000110101";
                        f_reg(206) <= "10101111101010000000010101010000";
                        f_reg(207) <= "10001100000111010000010110101100";
                        f_reg(208) <= "00011111101000000000000000000011";
                        f_reg(209) <= "00100000000111010000000000111100";
                        f_reg(210) <= "00010000000000000000000000000010";
                        f_reg(211) <= "00100000000111010000000000000000";
                        f_reg(212) <= "00010101001101110000000000101110";
                        f_reg(213) <= "10101111101010010000010101010100";
                        f_reg(214) <= "10001100000111010000010110101100";
                        f_reg(215) <= "00011111101000000000000000000011";
                        f_reg(216) <= "00100000000111010000000000111100";
                        f_reg(217) <= "00010000000000000000000000000010";
                        f_reg(218) <= "00100000000111010000000000000000";
                        f_reg(219) <= "00010101010110000000000000100111";
                        f_reg(220) <= "10101111101010100000010101011000";
                        f_reg(221) <= "10001100000111010000010110101100";
                        f_reg(222) <= "00011111101000000000000000000011";
                        f_reg(223) <= "00100000000111010000000000111100";
                        f_reg(224) <= "00010000000000000000000000000010";
                        f_reg(225) <= "00100000000111010000000000000000";
                        f_reg(226) <= "00010101011110010000000000100000";
                        f_reg(227) <= "10101111101010110000010101011100";
                        f_reg(228) <= "10001100000111010000010110101100";
                        f_reg(229) <= "00011111101000000000000000000011";
                        f_reg(230) <= "00100000000111010000000000111100";
                        f_reg(231) <= "00010000000000000000000000000010";
                        f_reg(232) <= "00100000000111010000000000000000";
                        f_reg(233) <= "00010101100110100000000000011001";
                        f_reg(234) <= "10101111101011000000010101100000";
                        f_reg(235) <= "10001100000111010000010110101100";
                        f_reg(236) <= "00011111101000000000000000000011";
                        f_reg(237) <= "00100000000111010000000000111100";
                        f_reg(238) <= "00010000000000000000000000000010";
                        f_reg(239) <= "00100000000111010000000000000000";
                        f_reg(240) <= "00010101101110110000000000010010";
                        f_reg(241) <= "10101111101011010000010101100100";
                        f_reg(242) <= "10001100000111010000010110101100";
                        f_reg(243) <= "00011111101000000000000000000011";
                        f_reg(244) <= "00100000000111010000000000111100";
                        f_reg(245) <= "00010000000000000000000000000010";
                        f_reg(246) <= "00100000000111010000000000000000";
                        f_reg(247) <= "00010101110111000000000000001011";
                        f_reg(248) <= "10101111101011100000010101101000";
                        f_reg(249) <= "10001100000111010000010110101100";
                        f_reg(250) <= "00011111101000000000000000000011";
                        f_reg(251) <= "00100000000111010000000000111100";
                        f_reg(252) <= "00010000000000000000000000000010";
                        f_reg(253) <= "00100000000111010000000000000000";
                        f_reg(254) <= "00010111110111110000000000000100";
                        f_reg(255) <= "10101111101111100000010101101100";
                        f_reg(256) <= "10101100000111010000010110101100";
                        f_reg(257) <= "00010000000000001111111110001010";
                        f_reg(258) <= "10001100000111010000010110101100";
                        f_reg(259) <= "10001111101000010000010100110100";
                        f_reg(260) <= "10001100000111010000010110101100";
                        f_reg(261) <= "10001111101011110000010100110100";
                        f_reg(262) <= "00010100001011111111111111111100";
                        f_reg(263) <= "10001100000111010000010110101100";
                        f_reg(264) <= "10001111101000100000010100111000";
                        f_reg(265) <= "10001100000111010000010110101100";
                        f_reg(266) <= "10001111101100000000010100111000";
                        f_reg(267) <= "00010100010100001111111111111100";
                        f_reg(268) <= "10001100000111010000010110101100";
                        f_reg(269) <= "10001111101000110000010100111100";
                        f_reg(270) <= "10001100000111010000010110101100";
                        f_reg(271) <= "10001111101100010000010100111100";
                        f_reg(272) <= "00010100011100011111111111111100";
                        f_reg(273) <= "10001100000111010000010110101100";
                        f_reg(274) <= "10001111101001000000010101000000";
                        f_reg(275) <= "10001100000111010000010110101100";
                        f_reg(276) <= "10001111101100100000010101000000";
                        f_reg(277) <= "00010100100100101111111111111100";
                        f_reg(278) <= "10001100000111010000010110101100";
                        f_reg(279) <= "10001111101001010000010101000100";
                        f_reg(280) <= "10001100000111010000010110101100";
                        f_reg(281) <= "10001111101100110000010101000100";
                        f_reg(282) <= "00010100101100111111111111111100";
                        f_reg(283) <= "10001100000111010000010110101100";
                        f_reg(284) <= "10001111101001100000010101001000";
                        f_reg(285) <= "10001100000111010000010110101100";
                        f_reg(286) <= "10001111101101000000010101001000";
                        f_reg(287) <= "00010100110101001111111111111100";
                        f_reg(288) <= "10001100000111010000010110101100";
                        f_reg(289) <= "10001111101001110000010101001100";
                        f_reg(290) <= "10001100000111010000010110101100";
                        f_reg(291) <= "10001111101101010000010101001100";
                        f_reg(292) <= "00010100111101011111111111111100";
                        f_reg(293) <= "10001100000111010000010110101100";
                        f_reg(294) <= "10001111101010000000010101010000";
                        f_reg(295) <= "10001100000111010000010110101100";
                        f_reg(296) <= "10001111101101100000010101010000";
                        f_reg(297) <= "00010101000101101111111111111100";
                        f_reg(298) <= "10001100000111010000010110101100";
                        f_reg(299) <= "10001111101010010000010101010100";
                        f_reg(300) <= "10001100000111010000010110101100";
                        f_reg(301) <= "10001111101101110000010101010100";
                        f_reg(302) <= "00010101001101111111111111111100";
                        f_reg(303) <= "10001100000111010000010110101100";
                        f_reg(304) <= "10001111101010100000010101011000";
                        f_reg(305) <= "10001100000111010000010110101100";
                        f_reg(306) <= "10001111101110000000010101011000";
                        f_reg(307) <= "00010101010110001111111111111100";
                        f_reg(308) <= "10001100000111010000010110101100";
                        f_reg(309) <= "10001111101010110000010101011100";
                        f_reg(310) <= "10001100000111010000010110101100";
                        f_reg(311) <= "10001111101110010000010101011100";
                        f_reg(312) <= "00010101011110011111111111111100";
                        f_reg(313) <= "10001100000111010000010110101100";
                        f_reg(314) <= "10001111101011000000010101100000";
                        f_reg(315) <= "10001100000111010000010110101100";
                        f_reg(316) <= "10001111101110100000010101100000";
                        f_reg(317) <= "00010101100110101111111111111100";
                        f_reg(318) <= "10001100000111010000010110101100";
                        f_reg(319) <= "10001111101011010000010101100100";
                        f_reg(320) <= "10001100000111010000010110101100";
                        f_reg(321) <= "10001111101110110000010101100100";
                        f_reg(322) <= "00010101101110111111111111111100";
                        f_reg(323) <= "10001100000111010000010110101100";
                        f_reg(324) <= "10001111101011100000010101101000";
                        f_reg(325) <= "10001100000111010000010110101100";
                        f_reg(326) <= "10001111101111000000010101101000";
                        f_reg(327) <= "00010101110111001111111111111100";
                        f_reg(328) <= "10001100000111010000010110101100";
                        f_reg(329) <= "10001111101111100000010101101100";
                        f_reg(330) <= "10001100000111010000010110101100";
                        f_reg(331) <= "10001111101111110000010101101100";
                        f_reg(332) <= "00010111110111111111111111111100";
                        f_reg(333) <= "00010000000000001111111100111110";
                        f_reg(334) <= "00000000000000000000000000000000";
                        f_reg(335) <= "00000000000000000000000000000000";
                        f_reg(336) <= "00000000000000000000000000000000";
                        f_reg(337) <= "00000000000000000000000000000000";
                        f_reg(338) <= "00000000000000000000000000000000";
                        f_reg(339) <= "00000000000000000000000000000000";
                        f_reg(340) <= "00000000000000000000000000000000";
                        f_reg(341) <= "00000000000000000000000000000000";
                        f_reg(342) <= "00000000000000000000000000000000";
                        f_reg(343) <= "00000000000000000000000000000000";
                        f_reg(344) <= "00000000000000000000000000000000";
                        f_reg(345) <= "00000000000000000000000000000000";
                        f_reg(346) <= "00000000000000000000000000000000";
                        f_reg(347) <= "00000000000000000000000000000000";
                        f_reg(348) <= "00000000000000000000000000000000";
                        f_reg(349) <= "00000000000000000000000000000000";
                        f_reg(350) <= "00000000000000000000000000000000";
                        f_reg(351) <= "00000000000000000000000000000000";
                        f_reg(352) <= "00000000000000000000000000000000";
                        f_reg(353) <= "00000000000000000000000000000000";
                        f_reg(354) <= "00000000000000000000000000000000";
                        f_reg(355) <= "00000000000000000000000000000000";
                        f_reg(356) <= "00000000000000000000000000000000";
                        f_reg(357) <= "00000000000000000000000000000000";
                        f_reg(358) <= "00000000000000000000000000000000";
                        f_reg(359) <= "00000000000000000000000000000000";
                        f_reg(360) <= "00000000000000000000000000000000";
                        f_reg(361) <= "00000000000000000000000000000000";
                        f_reg(362) <= "00000000000000000000000000000000";
                        f_reg(363) <= "00000000000000000000000000000000";
                        f_reg(364) <= "00000000000000000000001111100111";
                        f_reg(365) <= "00000000000000000000000000000000";
                        f_reg(366) <= "00000000000000000000000000000000";
                        f_reg(367) <= "00000000000000000000000000000000";
                        f_reg(368) <= "00000000000000000000000000000000";
                        f_reg(369) <= "00000000000000000000000000000000";
                        f_reg(370) <= "00000000000000000000000000000000";
                        f_reg(371) <= "00000000000000000000000000000000";
                        f_reg(372) <= "00000000000000000000000000000000";
                        f_reg(373) <= "00000000000000000000000000000000";
                        f_reg(374) <= "00000000000000000000000000000000";
                        f_reg(375) <= "00000000000000000000000000000000";
                        f_reg(376) <= "00000000000000000000000000000000";
                        f_reg(377) <= "00000000000000000000000000000000";
                        f_reg(378) <= "00000000000000000000000000000000";
                        f_reg(379) <= "00000000000000000000000000000000";
                        f_reg(380) <= "00000000000000000000000000000000";
                        f_reg(381) <= "00000000000000000000000000000000";
                        f_reg(382) <= "00000000000000000000000000000000";
                        f_reg(383) <= "00000000000000000000000000000000";
                        f_reg(384) <= "00000000000000000000000000000000";
                        f_reg(385) <= "00000000000000000000000000000000";
                        f_reg(386) <= "00000000000000000000000000000000";
                        f_reg(387) <= "00000000000000000000000000000000";
                        f_reg(388) <= "00000000000000000000000000000000";
                        f_reg(389) <= "00000000000000000000000000000000";
                        f_reg(390) <= "00000000000000000000000000000000";
                        f_reg(391) <= "00000000000000000000000000000000";
                        f_reg(392) <= "00000000000000000000000000000000";
                        f_reg(393) <= "00000000000000000000000000000000";
                        f_reg(394) <= "00000000000000000000000000000000";
                        f_reg(395) <= "00000000000000000000000000000000";
                        f_reg(396) <= "00000000000000000000000000000000";
                        f_reg(397) <= "00000000000000000000000000000000";
                        f_reg(398) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011101010000101101";
                        f_reg(4) <= "00000000000000000001010011000011";
                        f_reg(5) <= "00000000000000100001110111000000";
                        f_reg(6) <= "00111000001001000010001100100111";
                        f_reg(7) <= "00000000001001000010100000100101";
                        f_reg(8) <= "00111000010001100000110100110100";
                        f_reg(9) <= "00101100011001110100011001001000";
                        f_reg(10) <= "00100100110010001111010001101010";
                        f_reg(11) <= "00000000110001010100100000000110";
                        f_reg(12) <= "00100001000010101000111000000001";
                        f_reg(13) <= "00000000000001010101100000000111";
                        f_reg(14) <= "00000000110001100110000000000100";
                        f_reg(15) <= "00110101001011010100110100111001";
                        f_reg(16) <= "00000000000011000111000010000011";
                        f_reg(17) <= "10101100000000100000001000111100";
                        f_reg(18) <= "00110001110011110111100111000111";
                        f_reg(19) <= "00000000000000000000000000000000";
                        f_reg(20) <= "00000000000000000000000000000000";
                        f_reg(21) <= "00101001001100001101011001101000";
                        f_reg(22) <= "10101100000001110000001001000000";
                        f_reg(23) <= "00000000000010111000110111000010";
                        f_reg(24) <= "00100110001100101011010101001001";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00111100000100111000101011001111";
                        f_reg(27) <= "00000000000000000000000000000000";
                        f_reg(28) <= "00000000000100111010010101000010";
                        f_reg(29) <= "00000001101101001010100000100011";
                        f_reg(30) <= "00110100011101100011000000000110";
                        f_reg(31) <= "10101100000010100000001001000100";
                        f_reg(32) <= "00100110000101111111011111011000";
                        f_reg(33) <= "00000000000101111100000110000011";
                        f_reg(34) <= "00000000000000000000000000000000";
                        f_reg(35) <= "10101100000101100000001001001000";
                        f_reg(36) <= "00000010101110001100100000100111";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "10101100000011110000001001001100";
                        f_reg(39) <= "00000010010110011101000000101011";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "10101100000100010000001001010000";
                        f_reg(42) <= "00000000000000000000000000000000";
                        f_reg(43) <= "10101100000110100000001001010100";
                        f_reg(44) <= "00100011111111111111111111111111";
                        f_reg(45) <= "00011111111000001111111111010110";
                        f_reg(46) <= "00010000000000000000000101100001";
                        f_reg(47) <= "00111100000111100000001111100111";
                        f_reg(48) <= "00111100000111110000001111100111";
                        f_reg(49) <= "00000000000111101111010000000010";
                        f_reg(50) <= "00000000000111111111110000000010";
                        f_reg(51) <= "00111100000000011101010000101101";
                        f_reg(52) <= "00111100000011111101010000101101";
                        f_reg(53) <= "00000000000000000001010011000011";
                        f_reg(54) <= "00000000000000001000010011000011";
                        f_reg(55) <= "00000000000000100001110111000000";
                        f_reg(56) <= "00000000000100001000110111000000";
                        f_reg(57) <= "00111000001001000010001100100111";
                        f_reg(58) <= "00111001111100100010001100100111";
                        f_reg(59) <= "00000000001001000010100000100101";
                        f_reg(60) <= "00000001111100101001100000100101";
                        f_reg(61) <= "00111000010001100000110100110100";
                        f_reg(62) <= "00111010000101000000110100110100";
                        f_reg(63) <= "00101100011001110100011001001000";
                        f_reg(64) <= "00101110001101010100011001001000";
                        f_reg(65) <= "00100100110010001111010001101010";
                        f_reg(66) <= "00100110100101101111010001101010";
                        f_reg(67) <= "00000000110001010100100000000110";
                        f_reg(68) <= "00000010100100111011100000000110";
                        f_reg(69) <= "00100001000010101000111000000001";
                        f_reg(70) <= "00100010110110001000111000000001";
                        f_reg(71) <= "00000000000001010101100000000111";
                        f_reg(72) <= "00000000000100111100100000000111";
                        f_reg(73) <= "00000000110001100110000000000100";
                        f_reg(74) <= "00000010100101001101000000000100";
                        f_reg(75) <= "00110101001011010100110100111001";
                        f_reg(76) <= "00110110111110110100110100111001";
                        f_reg(77) <= "00000000000011000111000010000011";
                        f_reg(78) <= "00000000000110101110000010000011";
                        f_reg(79) <= "00010100010100000000000010110011";
                        f_reg(80) <= "10101100000000100000001000111100";
                        f_reg(81) <= "00110001110000010111100111000111";
                        f_reg(82) <= "00110011100011110111100111000111";
                        f_reg(83) <= "00000000000000000000000000000000";
                        f_reg(84) <= "00000000000000000000000000000000";
                        f_reg(85) <= "00000000000000000000000000000000";
                        f_reg(86) <= "00000000000000000000000000000000";
                        f_reg(87) <= "00101001001001001101011001101000";
                        f_reg(88) <= "00101010111100101101011001101000";
                        f_reg(89) <= "00010100111101010000000010101001";
                        f_reg(90) <= "10101100000001110000001001000000";
                        f_reg(91) <= "00000000000010110100010111000010";
                        f_reg(92) <= "00000000000110011011010111000010";
                        f_reg(93) <= "00100101000001011011010101001001";
                        f_reg(94) <= "00100110110100111011010101001001";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000000000000000000000000000";
                        f_reg(97) <= "00111100000001101000101011001111";
                        f_reg(98) <= "00111100000101001000101011001111";
                        f_reg(99) <= "00000000000000000000000000000000";
                        f_reg(100) <= "00000000000000000000000000000000";
                        f_reg(101) <= "00000000000001100110010101000010";
                        f_reg(102) <= "00000000000101001101010101000010";
                        f_reg(103) <= "00000001101011000001000000100011";
                        f_reg(104) <= "00000011011110101000000000100011";
                        f_reg(105) <= "00110100011011100011000000000110";
                        f_reg(106) <= "00110110001111000011000000000110";
                        f_reg(107) <= "00010101010110000000000010010111";
                        f_reg(108) <= "10101100000010100000001001000100";
                        f_reg(109) <= "00100100100010011111011111011000";
                        f_reg(110) <= "00100110010101111111011111011000";
                        f_reg(111) <= "00000000000010010011100110000011";
                        f_reg(112) <= "00000000000101111010100110000011";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00010101110111000000000010001111";
                        f_reg(116) <= "10101100000011100000001001001000";
                        f_reg(117) <= "00000000010001110101100000100111";
                        f_reg(118) <= "00000010000101011100100000100111";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000000000000000000000000000";
                        f_reg(121) <= "00010100001011110000000010001001";
                        f_reg(122) <= "10101100000000010000001001001100";
                        f_reg(123) <= "00000000101010110011000000101011";
                        f_reg(124) <= "00000010011110011010000000101011";
                        f_reg(125) <= "00000000000000000000000000000000";
                        f_reg(126) <= "00000000000000000000000000000000";
                        f_reg(127) <= "00010101000101100000000010000011";
                        f_reg(128) <= "10101100000010000000001001010000";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010100110101000000000001111111";
                        f_reg(132) <= "10101100000001100000001001010100";
                        f_reg(133) <= "00100011110111011111111100000110";
                        f_reg(134) <= "00010011101000000000000000010001";
                        f_reg(135) <= "00100011110111011111111000001100";
                        f_reg(136) <= "00010011101000000000000000001111";
                        f_reg(137) <= "00100011110111011111110100010010";
                        f_reg(138) <= "00010011101000000000000000001101";
                        f_reg(139) <= "00100011110111101111111111111111";
                        f_reg(140) <= "00100011111111111111111111111111";
                        f_reg(141) <= "00010111110111110000000001110101";
                        f_reg(142) <= "00011111111000001111111110100101";
                        f_reg(143) <= "00010000000000000000000100000000";
                        f_reg(144) <= "00000000000000000000000000000000";
                        f_reg(145) <= "00000000000000000000000000000000";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000000000000000000000000000";
                        f_reg(149) <= "00000000000000000000000000000000";
                        f_reg(150) <= "00000000000000000000000000000000";
                        f_reg(151) <= "10001100000111010000010110101100";
                        f_reg(152) <= "00011111101000000000000000000011";
                        f_reg(153) <= "00100000000111010000000000111100";
                        f_reg(154) <= "00010000000000000000000000000010";
                        f_reg(155) <= "00100000000111010000000000000000";
                        f_reg(156) <= "00010100001011110000000001100110";
                        f_reg(157) <= "10101111101000010000010100110100";
                        f_reg(158) <= "10001100000111010000010110101100";
                        f_reg(159) <= "00011111101000000000000000000011";
                        f_reg(160) <= "00100000000111010000000000111100";
                        f_reg(161) <= "00010000000000000000000000000010";
                        f_reg(162) <= "00100000000111010000000000000000";
                        f_reg(163) <= "00010100010100000000000001011111";
                        f_reg(164) <= "10101111101000100000010100111000";
                        f_reg(165) <= "10001100000111010000010110101100";
                        f_reg(166) <= "00011111101000000000000000000011";
                        f_reg(167) <= "00100000000111010000000000111100";
                        f_reg(168) <= "00010000000000000000000000000010";
                        f_reg(169) <= "00100000000111010000000000000000";
                        f_reg(170) <= "00010100011100010000000001011000";
                        f_reg(171) <= "10101111101000110000010100111100";
                        f_reg(172) <= "10001100000111010000010110101100";
                        f_reg(173) <= "00011111101000000000000000000011";
                        f_reg(174) <= "00100000000111010000000000111100";
                        f_reg(175) <= "00010000000000000000000000000010";
                        f_reg(176) <= "00100000000111010000000000000000";
                        f_reg(177) <= "00010100100100100000000001010001";
                        f_reg(178) <= "10101111101001000000010101000000";
                        f_reg(179) <= "10001100000111010000010110101100";
                        f_reg(180) <= "00011111101000000000000000000011";
                        f_reg(181) <= "00100000000111010000000000111100";
                        f_reg(182) <= "00010000000000000000000000000010";
                        f_reg(183) <= "00100000000111010000000000000000";
                        f_reg(184) <= "00010100101100110000000001001010";
                        f_reg(185) <= "10101111101001010000010101000100";
                        f_reg(186) <= "10001100000111010000010110101100";
                        f_reg(187) <= "00011111101000000000000000000011";
                        f_reg(188) <= "00100000000111010000000000111100";
                        f_reg(189) <= "00010000000000000000000000000010";
                        f_reg(190) <= "00100000000111010000000000000000";
                        f_reg(191) <= "00010100110101000000000001000011";
                        f_reg(192) <= "10101111101001100000010101001000";
                        f_reg(193) <= "10001100000111010000010110101100";
                        f_reg(194) <= "00011111101000000000000000000011";
                        f_reg(195) <= "00100000000111010000000000111100";
                        f_reg(196) <= "00010000000000000000000000000010";
                        f_reg(197) <= "00100000000111010000000000000000";
                        f_reg(198) <= "00010100111101010000000000111100";
                        f_reg(199) <= "10101111101001110000010101001100";
                        f_reg(200) <= "10001100000111010000010110101100";
                        f_reg(201) <= "00011111101000000000000000000011";
                        f_reg(202) <= "00100000000111010000000000111100";
                        f_reg(203) <= "00010000000000000000000000000010";
                        f_reg(204) <= "00100000000111010000000000000000";
                        f_reg(205) <= "00010101000101100000000000110101";
                        f_reg(206) <= "10101111101010000000010101010000";
                        f_reg(207) <= "10001100000111010000010110101100";
                        f_reg(208) <= "00011111101000000000000000000011";
                        f_reg(209) <= "00100000000111010000000000111100";
                        f_reg(210) <= "00010000000000000000000000000010";
                        f_reg(211) <= "00100000000111010000000000000000";
                        f_reg(212) <= "00010101001101110000000000101110";
                        f_reg(213) <= "10101111101010010000010101010100";
                        f_reg(214) <= "10001100000111010000010110101100";
                        f_reg(215) <= "00011111101000000000000000000011";
                        f_reg(216) <= "00100000000111010000000000111100";
                        f_reg(217) <= "00010000000000000000000000000010";
                        f_reg(218) <= "00100000000111010000000000000000";
                        f_reg(219) <= "00010101010110000000000000100111";
                        f_reg(220) <= "10101111101010100000010101011000";
                        f_reg(221) <= "10001100000111010000010110101100";
                        f_reg(222) <= "00011111101000000000000000000011";
                        f_reg(223) <= "00100000000111010000000000111100";
                        f_reg(224) <= "00010000000000000000000000000010";
                        f_reg(225) <= "00100000000111010000000000000000";
                        f_reg(226) <= "00010101011110010000000000100000";
                        f_reg(227) <= "10101111101010110000010101011100";
                        f_reg(228) <= "10001100000111010000010110101100";
                        f_reg(229) <= "00011111101000000000000000000011";
                        f_reg(230) <= "00100000000111010000000000111100";
                        f_reg(231) <= "00010000000000000000000000000010";
                        f_reg(232) <= "00100000000111010000000000000000";
                        f_reg(233) <= "00010101100110100000000000011001";
                        f_reg(234) <= "10101111101011000000010101100000";
                        f_reg(235) <= "10001100000111010000010110101100";
                        f_reg(236) <= "00011111101000000000000000000011";
                        f_reg(237) <= "00100000000111010000000000111100";
                        f_reg(238) <= "00010000000000000000000000000010";
                        f_reg(239) <= "00100000000111010000000000000000";
                        f_reg(240) <= "00010101101110110000000000010010";
                        f_reg(241) <= "10101111101011010000010101100100";
                        f_reg(242) <= "10001100000111010000010110101100";
                        f_reg(243) <= "00011111101000000000000000000011";
                        f_reg(244) <= "00100000000111010000000000111100";
                        f_reg(245) <= "00010000000000000000000000000010";
                        f_reg(246) <= "00100000000111010000000000000000";
                        f_reg(247) <= "00010101110111000000000000001011";
                        f_reg(248) <= "10101111101011100000010101101000";
                        f_reg(249) <= "10001100000111010000010110101100";
                        f_reg(250) <= "00011111101000000000000000000011";
                        f_reg(251) <= "00100000000111010000000000111100";
                        f_reg(252) <= "00010000000000000000000000000010";
                        f_reg(253) <= "00100000000111010000000000000000";
                        f_reg(254) <= "00010111110111110000000000000100";
                        f_reg(255) <= "10101111101111100000010101101100";
                        f_reg(256) <= "10101100000111010000010110101100";
                        f_reg(257) <= "00010000000000001111111110001010";
                        f_reg(258) <= "10001100000111010000010110101100";
                        f_reg(259) <= "10001111101000010000010100110100";
                        f_reg(260) <= "10001100000111010000010110101100";
                        f_reg(261) <= "10001111101011110000010100110100";
                        f_reg(262) <= "00010100001011111111111111111100";
                        f_reg(263) <= "10001100000111010000010110101100";
                        f_reg(264) <= "10001111101000100000010100111000";
                        f_reg(265) <= "10001100000111010000010110101100";
                        f_reg(266) <= "10001111101100000000010100111000";
                        f_reg(267) <= "00010100010100001111111111111100";
                        f_reg(268) <= "10001100000111010000010110101100";
                        f_reg(269) <= "10001111101000110000010100111100";
                        f_reg(270) <= "10001100000111010000010110101100";
                        f_reg(271) <= "10001111101100010000010100111100";
                        f_reg(272) <= "00010100011100011111111111111100";
                        f_reg(273) <= "10001100000111010000010110101100";
                        f_reg(274) <= "10001111101001000000010101000000";
                        f_reg(275) <= "10001100000111010000010110101100";
                        f_reg(276) <= "10001111101100100000010101000000";
                        f_reg(277) <= "00010100100100101111111111111100";
                        f_reg(278) <= "10001100000111010000010110101100";
                        f_reg(279) <= "10001111101001010000010101000100";
                        f_reg(280) <= "10001100000111010000010110101100";
                        f_reg(281) <= "10001111101100110000010101000100";
                        f_reg(282) <= "00010100101100111111111111111100";
                        f_reg(283) <= "10001100000111010000010110101100";
                        f_reg(284) <= "10001111101001100000010101001000";
                        f_reg(285) <= "10001100000111010000010110101100";
                        f_reg(286) <= "10001111101101000000010101001000";
                        f_reg(287) <= "00010100110101001111111111111100";
                        f_reg(288) <= "10001100000111010000010110101100";
                        f_reg(289) <= "10001111101001110000010101001100";
                        f_reg(290) <= "10001100000111010000010110101100";
                        f_reg(291) <= "10001111101101010000010101001100";
                        f_reg(292) <= "00010100111101011111111111111100";
                        f_reg(293) <= "10001100000111010000010110101100";
                        f_reg(294) <= "10001111101010000000010101010000";
                        f_reg(295) <= "10001100000111010000010110101100";
                        f_reg(296) <= "10001111101101100000010101010000";
                        f_reg(297) <= "00010101000101101111111111111100";
                        f_reg(298) <= "10001100000111010000010110101100";
                        f_reg(299) <= "10001111101010010000010101010100";
                        f_reg(300) <= "10001100000111010000010110101100";
                        f_reg(301) <= "10001111101101110000010101010100";
                        f_reg(302) <= "00010101001101111111111111111100";
                        f_reg(303) <= "10001100000111010000010110101100";
                        f_reg(304) <= "10001111101010100000010101011000";
                        f_reg(305) <= "10001100000111010000010110101100";
                        f_reg(306) <= "10001111101110000000010101011000";
                        f_reg(307) <= "00010101010110001111111111111100";
                        f_reg(308) <= "10001100000111010000010110101100";
                        f_reg(309) <= "10001111101010110000010101011100";
                        f_reg(310) <= "10001100000111010000010110101100";
                        f_reg(311) <= "10001111101110010000010101011100";
                        f_reg(312) <= "00010101011110011111111111111100";
                        f_reg(313) <= "10001100000111010000010110101100";
                        f_reg(314) <= "10001111101011000000010101100000";
                        f_reg(315) <= "10001100000111010000010110101100";
                        f_reg(316) <= "10001111101110100000010101100000";
                        f_reg(317) <= "00010101100110101111111111111100";
                        f_reg(318) <= "10001100000111010000010110101100";
                        f_reg(319) <= "10001111101011010000010101100100";
                        f_reg(320) <= "10001100000111010000010110101100";
                        f_reg(321) <= "10001111101110110000010101100100";
                        f_reg(322) <= "00010101101110111111111111111100";
                        f_reg(323) <= "10001100000111010000010110101100";
                        f_reg(324) <= "10001111101011100000010101101000";
                        f_reg(325) <= "10001100000111010000010110101100";
                        f_reg(326) <= "10001111101111000000010101101000";
                        f_reg(327) <= "00010101110111001111111111111100";
                        f_reg(328) <= "10001100000111010000010110101100";
                        f_reg(329) <= "10001111101111100000010101101100";
                        f_reg(330) <= "10001100000111010000010110101100";
                        f_reg(331) <= "10001111101111110000010101101100";
                        f_reg(332) <= "00010111110111111111111111111100";
                        f_reg(333) <= "00010000000000001111111100111110";
                        f_reg(334) <= "00000000000000000000000000000000";
                        f_reg(335) <= "00000000000000000000000000000000";
                        f_reg(336) <= "00000000000000000000000000000000";
                        f_reg(337) <= "00000000000000000000000000000000";
                        f_reg(338) <= "00000000000000000000000000000000";
                        f_reg(339) <= "00000000000000000000000000000000";
                        f_reg(340) <= "00000000000000000000000000000000";
                        f_reg(341) <= "00000000000000000000000000000000";
                        f_reg(342) <= "00000000000000000000000000000000";
                        f_reg(343) <= "00000000000000000000000000000000";
                        f_reg(344) <= "00000000000000000000000000000000";
                        f_reg(345) <= "00000000000000000000000000000000";
                        f_reg(346) <= "00000000000000000000000000000000";
                        f_reg(347) <= "00000000000000000000000000000000";
                        f_reg(348) <= "00000000000000000000000000000000";
                        f_reg(349) <= "00000000000000000000000000000000";
                        f_reg(350) <= "00000000000000000000000000000000";
                        f_reg(351) <= "00000000000000000000000000000000";
                        f_reg(352) <= "00000000000000000000000000000000";
                        f_reg(353) <= "00000000000000000000000000000000";
                        f_reg(354) <= "00000000000000000000000000000000";
                        f_reg(355) <= "00000000000000000000000000000000";
                        f_reg(356) <= "00000000000000000000000000000000";
                        f_reg(357) <= "00000000000000000000000000000000";
                        f_reg(358) <= "00000000000000000000000000000000";
                        f_reg(359) <= "00000000000000000000000000000000";
                        f_reg(360) <= "00000000000000000000000000000000";
                        f_reg(361) <= "00000000000000000000000000000000";
                        f_reg(362) <= "00000000000000000000000000000000";
                        f_reg(363) <= "00000000000000000000000000000000";
                        f_reg(364) <= "00000000000000000000001111100111";
                        f_reg(365) <= "00000000000000000000000000000000";
                        f_reg(366) <= "00000000000000000000000000000000";
                        f_reg(367) <= "00000000000000000000000000000000";
                        f_reg(368) <= "00000000000000000000000000000000";
                        f_reg(369) <= "00000000000000000000000000000000";
                        f_reg(370) <= "00000000000000000000000000000000";
                        f_reg(371) <= "00000000000000000000000000000000";
                        f_reg(372) <= "00000000000000000000000000000000";
                        f_reg(373) <= "00000000000000000000000000000000";
                        f_reg(374) <= "00000000000000000000000000000000";
                        f_reg(375) <= "00000000000000000000000000000000";
                        f_reg(376) <= "00000000000000000000000000000000";
                        f_reg(377) <= "00000000000000000000000000000000";
                        f_reg(378) <= "00000000000000000000000000000000";
                        f_reg(379) <= "00000000000000000000000000000000";
                        f_reg(380) <= "00000000000000000000000000000000";
                        f_reg(381) <= "00000000000000000000000000000000";
                        f_reg(382) <= "00000000000000000000000000000000";
                        f_reg(383) <= "00000000000000000000000000000000";
                        f_reg(384) <= "00000000000000000000000000000000";
                        f_reg(385) <= "00000000000000000000000000000000";
                        f_reg(386) <= "00000000000000000000000000000000";
                        f_reg(387) <= "00000000000000000000000000000000";
                        f_reg(388) <= "00000000000000000000000000000000";
                        f_reg(389) <= "00000000000000000000000000000000";
                        f_reg(390) <= "00000000000000000000000000000000";
                        f_reg(391) <= "00000000000000000000000000000000";
                        f_reg(392) <= "00000000000000000000000000000000";
                        f_reg(393) <= "00000000000000000000000000000000";
                        f_reg(394) <= "00000000000000000000000000000000";
                        f_reg(395) <= "00000000000000000000000000000000";
                        f_reg(396) <= "00000000000000000000000000000000";
                        f_reg(397) <= "00000000000000000000000000000000";
                        f_reg(398) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 -11219
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SRA R2 R0 19
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SLL R3 R2 23
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- XORI R4 R1 8999
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- OR R5 R1 R4
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- XORI R6 R2 3380
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- SLTIU R7 R3 17992
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- ADDIU R8 R6 -2966
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- SRLV R9 R5 R6
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- ADDI R10 R8 -29183
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- SRAV R11 R5 R0
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- SLLV R12 R6 R6
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- ORI R13 R9 19769
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- SRA R14 R12 2
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- SW R2 R0 572
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- ANDI R15 R14 31175
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- NOP
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- NOP
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SLTI R16 R9 -10648
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- SW R7 R0 576
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- SRL R17 R11 23
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- ADDIU R18 R17 -19127
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- NOP
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- LUI R19 -30001
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- NOP
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- SRL R20 R19 21
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- SUBU R21 R13 R20
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- ORI R22 R3 12294
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- SW R10 R0 580
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- ADDIU R23 R16 -2088
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- SRA R24 R23 6
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- NOP
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- SW R22 R0 584
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- NOR R25 R21 R24
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- NOP
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- SW R15 R0 588
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- SLTU R26 R18 R25
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- NOP
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- SW R17 R0 592
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- NOP
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SW R26 R0 596
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- ADDI R31 R31 -1
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- BGTZ R31 -42
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- BEQ R0 R0 353
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- LUI R30 999
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- LUI R31 999
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- SRL R30 R30 16
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- SRL R31 R31 16
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- LUI R1 -11219
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- LUI R15 -11219
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- SRA R2 R0 19
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SRA R16 R0 19
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SLL R3 R2 23
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- SLL R17 R16 23
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- XORI R4 R1 8999
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- XORI R18 R15 8999
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- OR R5 R1 R4
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- OR R19 R15 R18
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- XORI R6 R2 3380
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- XORI R20 R16 3380
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- SLTIU R7 R3 17992
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- SLTIU R21 R17 17992
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- ADDIU R8 R6 -2966
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- ADDIU R22 R20 -2966
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- SRLV R9 R5 R6
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- SRLV R23 R19 R20
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- ADDI R10 R8 -29183
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- ADDI R24 R22 -29183
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- SRAV R11 R5 R0
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- SRAV R25 R19 R0
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SLLV R12 R6 R6
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- SLLV R26 R20 R20
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- ORI R13 R9 19769
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- ORI R27 R23 19769
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- SRA R14 R12 2
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- SRA R28 R26 2
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- BNE R2 R16 179
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- SW R2 R0 572
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- ANDI R1 R14 31175
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- ANDI R15 R28 31175
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- NOP
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- NOP
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- NOP
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- NOP
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SLTI R4 R9 -10648
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- SLTI R18 R23 -10648
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- BNE R7 R21 169
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- SW R7 R0 576
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- SRL R8 R11 23
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- SRL R22 R25 23
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- ADDIU R5 R8 -19127
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- ADDIU R19 R22 -19127
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- NOP
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- NOP
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- LUI R6 -30001
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- LUI R20 -30001
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- NOP
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- NOP
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- SRL R12 R6 21
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- SRL R26 R20 21
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SUBU R2 R13 R12
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- SUBU R16 R27 R26
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- ORI R14 R3 12294
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- ORI R28 R17 12294
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- BNE R10 R24 151
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- SW R10 R0 580
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- ADDIU R9 R4 -2088
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- ADDIU R23 R18 -2088
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- SRA R7 R9 6
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- SRA R21 R23 6
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- NOP
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- NOP
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- BNE R14 R28 143
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- SW R14 R0 584
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- NOR R11 R2 R7
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- NOR R25 R16 R21
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- NOP
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- NOP
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- BNE R1 R15 137
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- SW R1 R0 588
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- SLTU R6 R5 R11
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SLTU R20 R19 R25
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- NOP
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- NOP
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- BNE R8 R22 131
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SW R8 R0 592
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- NOP
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- NOP
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- BNE R6 R20 127
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- SW R6 R0 596
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- ADDI R29 R30 -250
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- BEQ R29 R0 17
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- ADDI R29 R30 -500
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- BEQ R29 R0 15
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- ADDI R29 R30 -750
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- BEQ R29 R0 13
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- ADDI R30 R30 -1
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- ADDI R31 R31 -1
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- BNE R30 R31 117
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- BGTZ R31 -91
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- BEQ R0 R0 256
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- NOP
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- NOP
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- NOP
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- NOP
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- NOP
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- NOP
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- NOP
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- LW R29 R0 1452
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- BGTZ R29 3
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- ADDI R29 R0 60
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- BEQ R0 R0 2
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- ADDI R29 R0 0
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- BNE R1 R15 102
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- SW R1 R29 1332
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- LW R29 R0 1452
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- BGTZ R29 3
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- ADDI R29 R0 60
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- BEQ R0 R0 2
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- ADDI R29 R0 0
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- BNE R2 R16 95
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- SW R2 R29 1336
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- LW R29 R0 1452
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- BGTZ R29 3
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- ADDI R29 R0 60
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- BEQ R0 R0 2
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- ADDI R29 R0 0
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- BNE R3 R17 88
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- SW R3 R29 1340
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- LW R29 R0 1452
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- BGTZ R29 3
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- ADDI R29 R0 60
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- BEQ R0 R0 2
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- ADDI R29 R0 0
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- BNE R4 R18 81
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- SW R4 R29 1344
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- LW R29 R0 1452
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- BGTZ R29 3
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- ADDI R29 R0 60
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- BEQ R0 R0 2
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- ADDI R29 R0 0
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- BNE R5 R19 74
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- SW R5 R29 1348
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- LW R29 R0 1452
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- BGTZ R29 3
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- ADDI R29 R0 60
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- BEQ R0 R0 2
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- ADDI R29 R0 0
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- BNE R6 R20 67
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- SW R6 R29 1352
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- LW R29 R0 1452
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- BGTZ R29 3
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- ADDI R29 R0 60
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- BEQ R0 R0 2
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- ADDI R29 R0 0
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- BNE R7 R21 60
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- SW R7 R29 1356
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- LW R29 R0 1452
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- BGTZ R29 3
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- ADDI R29 R0 60
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- BEQ R0 R0 2
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- ADDI R29 R0 0
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- BNE R8 R22 53
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- SW R8 R29 1360
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- LW R29 R0 1452
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- BGTZ R29 3
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- ADDI R29 R0 60
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- BEQ R0 R0 2
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- ADDI R29 R0 0
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- BNE R9 R23 46
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- SW R9 R29 1364
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- LW R29 R0 1452
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- BGTZ R29 3
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- ADDI R29 R0 60
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- BEQ R0 R0 2
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- ADDI R29 R0 0
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- BNE R10 R24 39
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- SW R10 R29 1368
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- LW R29 R0 1452
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- BGTZ R29 3
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- ADDI R29 R0 60
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- BEQ R0 R0 2
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- ADDI R29 R0 0
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- BNE R11 R25 32
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- SW R11 R29 1372
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- LW R29 R0 1452
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- BGTZ R29 3
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- ADDI R29 R0 60
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- BEQ R0 R0 2
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- ADDI R29 R0 0
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- BNE R12 R26 25
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- SW R12 R29 1376
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- LW R29 R0 1452
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- BGTZ R29 3
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- ADDI R29 R0 60
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- BEQ R0 R0 2
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- ADDI R29 R0 0
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- BNE R13 R27 18
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- SW R13 R29 1380
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- LW R29 R0 1452
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- BGTZ R29 3
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- ADDI R29 R0 60
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- BEQ R0 R0 2
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- ADDI R29 R0 0
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- BNE R14 R28 11
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- SW R14 R29 1384
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- LW R29 R0 1452
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- BGTZ R29 3
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- ADDI R29 R0 60
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- BEQ R0 R0 2
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- ADDI R29 R0 0
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- BNE R30 R31 4
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- SW R30 R29 1388
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- SW R29 R0 1452
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- BEQ R0 R0 -118
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- LW R29 R0 1452
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- LW R1 R29 1332
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- LW R29 R0 1452
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- LW R15 R29 1332
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- BNE R1 R15 -4
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- LW R29 R0 1452
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- LW R2 R29 1336
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- LW R29 R0 1452
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- LW R16 R29 1336
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- BNE R2 R16 -4
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- LW R29 R0 1452
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- LW R3 R29 1340
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- LW R29 R0 1452
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- LW R17 R29 1340
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- BNE R3 R17 -4
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- LW R29 R0 1452
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- LW R4 R29 1344
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- LW R29 R0 1452
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- LW R18 R29 1344
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- BNE R4 R18 -4
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- LW R29 R0 1452
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- LW R5 R29 1348
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- LW R29 R0 1452
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- LW R19 R29 1348
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- BNE R5 R19 -4
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- LW R29 R0 1452
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- LW R6 R29 1352
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- LW R29 R0 1452
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- LW R20 R29 1352
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- BNE R6 R20 -4
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- LW R29 R0 1452
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- LW R7 R29 1356
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- LW R29 R0 1452
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- LW R21 R29 1356
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- BNE R7 R21 -4
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- LW R29 R0 1452
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- LW R8 R29 1360
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- LW R29 R0 1452
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- LW R22 R29 1360
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- BNE R8 R22 -4
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- LW R29 R0 1452
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- LW R9 R29 1364
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- LW R29 R0 1452
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- LW R23 R29 1364
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- BNE R9 R23 -4
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- LW R29 R0 1452
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- LW R10 R29 1368
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- LW R29 R0 1452
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- LW R24 R29 1368
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- BNE R10 R24 -4
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- LW R29 R0 1452
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- LW R11 R29 1372
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- LW R29 R0 1452
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- LW R25 R29 1372
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- BNE R11 R25 -4
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- LW R29 R0 1452
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- LW R12 R29 1376
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- LW R29 R0 1452
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- LW R26 R29 1376
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- BNE R12 R26 -4
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- LW R29 R0 1452
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- LW R13 R29 1380
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- LW R29 R0 1452
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- LW R27 R29 1380
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- BNE R13 R27 -4
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- LW R29 R0 1452
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- LW R14 R29 1384
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- LW R29 R0 1452
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- LW R28 R29 1384
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- BNE R14 R28 -4
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- LW R29 R0 1452
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- LW R30 R29 1388
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- LW R29 R0 1452
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- LW R31 R29 1388
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- BNE R30 R31 -4
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- BEQ R0 R0 -194
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- NOP
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- NOP
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- NOP
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- NOP
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- NOP
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- NOP
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- NOP
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- NOP
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- NOP
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- NOP
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- NOP
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- NOP
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- NOP
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- NOP
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- NOP
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- NOP
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- NOP
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- NOP
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- NOP
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- NOP
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- NOP
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- NOP
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- NOP
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- NOP
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- NOP
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- NOP
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- NOP
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- NOP
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- NOP
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- NOP
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- NOP
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- NOP
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- NOP
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- NOP
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- NOP
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- NOP
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- NOP
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- NOP
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- NOP
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- NOP
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- NOP
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- NOP
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- NOP
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- NOP
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- NOP
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- NOP
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- NOP
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- NOP
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- NOP
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- NOP
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- NOP
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- NOP
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- NOP
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- NOP
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- NOP
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- NOP
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- NOP
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- NOP
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- NOP
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- NOP
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- NOP
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- NOP
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- NOP
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- NOP
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- NOP
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011101010000101101";
                        f_reg(4) <= "00000000000000000001010011000011";
                        f_reg(5) <= "00000000000000100001110111000000";
                        f_reg(6) <= "00111000001001000010001100100111";
                        f_reg(7) <= "00000000001001000010100000100101";
                        f_reg(8) <= "00111000010001100000110100110100";
                        f_reg(9) <= "00101100011001110100011001001000";
                        f_reg(10) <= "00100100110010001111010001101010";
                        f_reg(11) <= "00000000110001010100100000000110";
                        f_reg(12) <= "00100001000010101000111000000001";
                        f_reg(13) <= "00000000000001010101100000000111";
                        f_reg(14) <= "00000000110001100110000000000100";
                        f_reg(15) <= "00110101001011010100110100111001";
                        f_reg(16) <= "00000000000011000111000010000011";
                        f_reg(17) <= "10101100000000100000001000111100";
                        f_reg(18) <= "00110001110011110111100111000111";
                        f_reg(19) <= "00000000000000000000000000000000";
                        f_reg(20) <= "00000000000000000000000000000000";
                        f_reg(21) <= "00101001001100001101011001101000";
                        f_reg(22) <= "10101100000001110000001001000000";
                        f_reg(23) <= "00000000000010111000110111000010";
                        f_reg(24) <= "00100110001100101011010101001001";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00111100000100111000101011001111";
                        f_reg(27) <= "00000000000000000000000000000000";
                        f_reg(28) <= "00000000000100111010010101000010";
                        f_reg(29) <= "00000001101101001010100000100011";
                        f_reg(30) <= "00110100011101100011000000000110";
                        f_reg(31) <= "10101100000010100000001001000100";
                        f_reg(32) <= "00100110000101111111011111011000";
                        f_reg(33) <= "00000000000101111100000110000011";
                        f_reg(34) <= "00000000000000000000000000000000";
                        f_reg(35) <= "10101100000101100000001001001000";
                        f_reg(36) <= "00000010101110001100100000100111";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "10101100000011110000001001001100";
                        f_reg(39) <= "00000010010110011101000000101011";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "10101100000100010000001001010000";
                        f_reg(42) <= "00000000000000000000000000000000";
                        f_reg(43) <= "10101100000110100000001001010100";
                        f_reg(44) <= "00100011111111111111111111111111";
                        f_reg(45) <= "00011111111000001111111111010110";
                        f_reg(46) <= "00010000000000000000000101100001";
                        f_reg(47) <= "00111100000111100000001111100111";
                        f_reg(48) <= "00111100000111110000001111100111";
                        f_reg(49) <= "00000000000111101111010000000010";
                        f_reg(50) <= "00000000000111111111110000000010";
                        f_reg(51) <= "00111100000000011101010000101101";
                        f_reg(52) <= "00111100000011111101010000101101";
                        f_reg(53) <= "00000000000000000001010011000011";
                        f_reg(54) <= "00000000000000001000010011000011";
                        f_reg(55) <= "00000000000000100001110111000000";
                        f_reg(56) <= "00000000000100001000110111000000";
                        f_reg(57) <= "00111000001001000010001100100111";
                        f_reg(58) <= "00111001111100100010001100100111";
                        f_reg(59) <= "00000000001001000010100000100101";
                        f_reg(60) <= "00000001111100101001100000100101";
                        f_reg(61) <= "00111000010001100000110100110100";
                        f_reg(62) <= "00111010000101000000110100110100";
                        f_reg(63) <= "00101100011001110100011001001000";
                        f_reg(64) <= "00101110001101010100011001001000";
                        f_reg(65) <= "00100100110010001111010001101010";
                        f_reg(66) <= "00100110100101101111010001101010";
                        f_reg(67) <= "00000000110001010100100000000110";
                        f_reg(68) <= "00000010100100111011100000000110";
                        f_reg(69) <= "00100001000010101000111000000001";
                        f_reg(70) <= "00100010110110001000111000000001";
                        f_reg(71) <= "00000000000001010101100000000111";
                        f_reg(72) <= "00000000000100111100100000000111";
                        f_reg(73) <= "00000000110001100110000000000100";
                        f_reg(74) <= "00000010100101001101000000000100";
                        f_reg(75) <= "00110101001011010100110100111001";
                        f_reg(76) <= "00110110111110110100110100111001";
                        f_reg(77) <= "00000000000011000111000010000011";
                        f_reg(78) <= "00000000000110101110000010000011";
                        f_reg(79) <= "00010100010100000000000010110011";
                        f_reg(80) <= "10101100000000100000001000111100";
                        f_reg(81) <= "00110001110000010111100111000111";
                        f_reg(82) <= "00110011100011110111100111000111";
                        f_reg(83) <= "00000000000000000000000000000000";
                        f_reg(84) <= "00000000000000000000000000000000";
                        f_reg(85) <= "00000000000000000000000000000000";
                        f_reg(86) <= "00000000000000000000000000000000";
                        f_reg(87) <= "00101001001001001101011001101000";
                        f_reg(88) <= "00101010111100101101011001101000";
                        f_reg(89) <= "00010100111101010000000010101001";
                        f_reg(90) <= "10101100000001110000001001000000";
                        f_reg(91) <= "00000000000010110100010111000010";
                        f_reg(92) <= "00000000000110011011010111000010";
                        f_reg(93) <= "00100101000001011011010101001001";
                        f_reg(94) <= "00100110110100111011010101001001";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000000000000000000000000000";
                        f_reg(97) <= "00111100000001101000101011001111";
                        f_reg(98) <= "00111100000101001000101011001111";
                        f_reg(99) <= "00000000000000000000000000000000";
                        f_reg(100) <= "00000000000000000000000000000000";
                        f_reg(101) <= "00000000000001100110010101000010";
                        f_reg(102) <= "00000000000101001101010101000010";
                        f_reg(103) <= "00000001101011000001000000100011";
                        f_reg(104) <= "00000011011110101000000000100011";
                        f_reg(105) <= "00110100011011100011000000000110";
                        f_reg(106) <= "00110110001111000011000000000110";
                        f_reg(107) <= "00010101010110000000000010010111";
                        f_reg(108) <= "10101100000010100000001001000100";
                        f_reg(109) <= "00100100100010011111011111011000";
                        f_reg(110) <= "00100110010101111111011111011000";
                        f_reg(111) <= "00000000000010010011100110000011";
                        f_reg(112) <= "00000000000101111010100110000011";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00010101110111000000000010001111";
                        f_reg(116) <= "10101100000011100000001001001000";
                        f_reg(117) <= "00000000010001110101100000100111";
                        f_reg(118) <= "00000010000101011100100000100111";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000000000000000000000000000";
                        f_reg(121) <= "00010100001011110000000010001001";
                        f_reg(122) <= "10101100000000010000001001001100";
                        f_reg(123) <= "00000000101010110011000000101011";
                        f_reg(124) <= "00000010011110011010000000101011";
                        f_reg(125) <= "00000000000000000000000000000000";
                        f_reg(126) <= "00000000000000000000000000000000";
                        f_reg(127) <= "00010101000101100000000010000011";
                        f_reg(128) <= "10101100000010000000001001010000";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010100110101000000000001111111";
                        f_reg(132) <= "10101100000001100000001001010100";
                        f_reg(133) <= "00100011110111011111111100000110";
                        f_reg(134) <= "00010011101000000000000000010001";
                        f_reg(135) <= "00100011110111011111111000001100";
                        f_reg(136) <= "00010011101000000000000000001111";
                        f_reg(137) <= "00100011110111011111110100010010";
                        f_reg(138) <= "00010011101000000000000000001101";
                        f_reg(139) <= "00100011110111101111111111111111";
                        f_reg(140) <= "00100011111111111111111111111111";
                        f_reg(141) <= "00010111110111110000000001110101";
                        f_reg(142) <= "00011111111000001111111110100101";
                        f_reg(143) <= "00010000000000000000000100000000";
                        f_reg(144) <= "00000000000000000000000000000000";
                        f_reg(145) <= "00000000000000000000000000000000";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000000000000000000000000000";
                        f_reg(149) <= "00000000000000000000000000000000";
                        f_reg(150) <= "00000000000000000000000000000000";
                        f_reg(151) <= "10001100000111010000010110101100";
                        f_reg(152) <= "00011111101000000000000000000011";
                        f_reg(153) <= "00100000000111010000000000111100";
                        f_reg(154) <= "00010000000000000000000000000010";
                        f_reg(155) <= "00100000000111010000000000000000";
                        f_reg(156) <= "00010100001011110000000001100110";
                        f_reg(157) <= "10101111101000010000010100110100";
                        f_reg(158) <= "10001100000111010000010110101100";
                        f_reg(159) <= "00011111101000000000000000000011";
                        f_reg(160) <= "00100000000111010000000000111100";
                        f_reg(161) <= "00010000000000000000000000000010";
                        f_reg(162) <= "00100000000111010000000000000000";
                        f_reg(163) <= "00010100010100000000000001011111";
                        f_reg(164) <= "10101111101000100000010100111000";
                        f_reg(165) <= "10001100000111010000010110101100";
                        f_reg(166) <= "00011111101000000000000000000011";
                        f_reg(167) <= "00100000000111010000000000111100";
                        f_reg(168) <= "00010000000000000000000000000010";
                        f_reg(169) <= "00100000000111010000000000000000";
                        f_reg(170) <= "00010100011100010000000001011000";
                        f_reg(171) <= "10101111101000110000010100111100";
                        f_reg(172) <= "10001100000111010000010110101100";
                        f_reg(173) <= "00011111101000000000000000000011";
                        f_reg(174) <= "00100000000111010000000000111100";
                        f_reg(175) <= "00010000000000000000000000000010";
                        f_reg(176) <= "00100000000111010000000000000000";
                        f_reg(177) <= "00010100100100100000000001010001";
                        f_reg(178) <= "10101111101001000000010101000000";
                        f_reg(179) <= "10001100000111010000010110101100";
                        f_reg(180) <= "00011111101000000000000000000011";
                        f_reg(181) <= "00100000000111010000000000111100";
                        f_reg(182) <= "00010000000000000000000000000010";
                        f_reg(183) <= "00100000000111010000000000000000";
                        f_reg(184) <= "00010100101100110000000001001010";
                        f_reg(185) <= "10101111101001010000010101000100";
                        f_reg(186) <= "10001100000111010000010110101100";
                        f_reg(187) <= "00011111101000000000000000000011";
                        f_reg(188) <= "00100000000111010000000000111100";
                        f_reg(189) <= "00010000000000000000000000000010";
                        f_reg(190) <= "00100000000111010000000000000000";
                        f_reg(191) <= "00010100110101000000000001000011";
                        f_reg(192) <= "10101111101001100000010101001000";
                        f_reg(193) <= "10001100000111010000010110101100";
                        f_reg(194) <= "00011111101000000000000000000011";
                        f_reg(195) <= "00100000000111010000000000111100";
                        f_reg(196) <= "00010000000000000000000000000010";
                        f_reg(197) <= "00100000000111010000000000000000";
                        f_reg(198) <= "00010100111101010000000000111100";
                        f_reg(199) <= "10101111101001110000010101001100";
                        f_reg(200) <= "10001100000111010000010110101100";
                        f_reg(201) <= "00011111101000000000000000000011";
                        f_reg(202) <= "00100000000111010000000000111100";
                        f_reg(203) <= "00010000000000000000000000000010";
                        f_reg(204) <= "00100000000111010000000000000000";
                        f_reg(205) <= "00010101000101100000000000110101";
                        f_reg(206) <= "10101111101010000000010101010000";
                        f_reg(207) <= "10001100000111010000010110101100";
                        f_reg(208) <= "00011111101000000000000000000011";
                        f_reg(209) <= "00100000000111010000000000111100";
                        f_reg(210) <= "00010000000000000000000000000010";
                        f_reg(211) <= "00100000000111010000000000000000";
                        f_reg(212) <= "00010101001101110000000000101110";
                        f_reg(213) <= "10101111101010010000010101010100";
                        f_reg(214) <= "10001100000111010000010110101100";
                        f_reg(215) <= "00011111101000000000000000000011";
                        f_reg(216) <= "00100000000111010000000000111100";
                        f_reg(217) <= "00010000000000000000000000000010";
                        f_reg(218) <= "00100000000111010000000000000000";
                        f_reg(219) <= "00010101010110000000000000100111";
                        f_reg(220) <= "10101111101010100000010101011000";
                        f_reg(221) <= "10001100000111010000010110101100";
                        f_reg(222) <= "00011111101000000000000000000011";
                        f_reg(223) <= "00100000000111010000000000111100";
                        f_reg(224) <= "00010000000000000000000000000010";
                        f_reg(225) <= "00100000000111010000000000000000";
                        f_reg(226) <= "00010101011110010000000000100000";
                        f_reg(227) <= "10101111101010110000010101011100";
                        f_reg(228) <= "10001100000111010000010110101100";
                        f_reg(229) <= "00011111101000000000000000000011";
                        f_reg(230) <= "00100000000111010000000000111100";
                        f_reg(231) <= "00010000000000000000000000000010";
                        f_reg(232) <= "00100000000111010000000000000000";
                        f_reg(233) <= "00010101100110100000000000011001";
                        f_reg(234) <= "10101111101011000000010101100000";
                        f_reg(235) <= "10001100000111010000010110101100";
                        f_reg(236) <= "00011111101000000000000000000011";
                        f_reg(237) <= "00100000000111010000000000111100";
                        f_reg(238) <= "00010000000000000000000000000010";
                        f_reg(239) <= "00100000000111010000000000000000";
                        f_reg(240) <= "00010101101110110000000000010010";
                        f_reg(241) <= "10101111101011010000010101100100";
                        f_reg(242) <= "10001100000111010000010110101100";
                        f_reg(243) <= "00011111101000000000000000000011";
                        f_reg(244) <= "00100000000111010000000000111100";
                        f_reg(245) <= "00010000000000000000000000000010";
                        f_reg(246) <= "00100000000111010000000000000000";
                        f_reg(247) <= "00010101110111000000000000001011";
                        f_reg(248) <= "10101111101011100000010101101000";
                        f_reg(249) <= "10001100000111010000010110101100";
                        f_reg(250) <= "00011111101000000000000000000011";
                        f_reg(251) <= "00100000000111010000000000111100";
                        f_reg(252) <= "00010000000000000000000000000010";
                        f_reg(253) <= "00100000000111010000000000000000";
                        f_reg(254) <= "00010111110111110000000000000100";
                        f_reg(255) <= "10101111101111100000010101101100";
                        f_reg(256) <= "10101100000111010000010110101100";
                        f_reg(257) <= "00010000000000001111111110001010";
                        f_reg(258) <= "10001100000111010000010110101100";
                        f_reg(259) <= "10001111101000010000010100110100";
                        f_reg(260) <= "10001100000111010000010110101100";
                        f_reg(261) <= "10001111101011110000010100110100";
                        f_reg(262) <= "00010100001011111111111111111100";
                        f_reg(263) <= "10001100000111010000010110101100";
                        f_reg(264) <= "10001111101000100000010100111000";
                        f_reg(265) <= "10001100000111010000010110101100";
                        f_reg(266) <= "10001111101100000000010100111000";
                        f_reg(267) <= "00010100010100001111111111111100";
                        f_reg(268) <= "10001100000111010000010110101100";
                        f_reg(269) <= "10001111101000110000010100111100";
                        f_reg(270) <= "10001100000111010000010110101100";
                        f_reg(271) <= "10001111101100010000010100111100";
                        f_reg(272) <= "00010100011100011111111111111100";
                        f_reg(273) <= "10001100000111010000010110101100";
                        f_reg(274) <= "10001111101001000000010101000000";
                        f_reg(275) <= "10001100000111010000010110101100";
                        f_reg(276) <= "10001111101100100000010101000000";
                        f_reg(277) <= "00010100100100101111111111111100";
                        f_reg(278) <= "10001100000111010000010110101100";
                        f_reg(279) <= "10001111101001010000010101000100";
                        f_reg(280) <= "10001100000111010000010110101100";
                        f_reg(281) <= "10001111101100110000010101000100";
                        f_reg(282) <= "00010100101100111111111111111100";
                        f_reg(283) <= "10001100000111010000010110101100";
                        f_reg(284) <= "10001111101001100000010101001000";
                        f_reg(285) <= "10001100000111010000010110101100";
                        f_reg(286) <= "10001111101101000000010101001000";
                        f_reg(287) <= "00010100110101001111111111111100";
                        f_reg(288) <= "10001100000111010000010110101100";
                        f_reg(289) <= "10001111101001110000010101001100";
                        f_reg(290) <= "10001100000111010000010110101100";
                        f_reg(291) <= "10001111101101010000010101001100";
                        f_reg(292) <= "00010100111101011111111111111100";
                        f_reg(293) <= "10001100000111010000010110101100";
                        f_reg(294) <= "10001111101010000000010101010000";
                        f_reg(295) <= "10001100000111010000010110101100";
                        f_reg(296) <= "10001111101101100000010101010000";
                        f_reg(297) <= "00010101000101101111111111111100";
                        f_reg(298) <= "10001100000111010000010110101100";
                        f_reg(299) <= "10001111101010010000010101010100";
                        f_reg(300) <= "10001100000111010000010110101100";
                        f_reg(301) <= "10001111101101110000010101010100";
                        f_reg(302) <= "00010101001101111111111111111100";
                        f_reg(303) <= "10001100000111010000010110101100";
                        f_reg(304) <= "10001111101010100000010101011000";
                        f_reg(305) <= "10001100000111010000010110101100";
                        f_reg(306) <= "10001111101110000000010101011000";
                        f_reg(307) <= "00010101010110001111111111111100";
                        f_reg(308) <= "10001100000111010000010110101100";
                        f_reg(309) <= "10001111101010110000010101011100";
                        f_reg(310) <= "10001100000111010000010110101100";
                        f_reg(311) <= "10001111101110010000010101011100";
                        f_reg(312) <= "00010101011110011111111111111100";
                        f_reg(313) <= "10001100000111010000010110101100";
                        f_reg(314) <= "10001111101011000000010101100000";
                        f_reg(315) <= "10001100000111010000010110101100";
                        f_reg(316) <= "10001111101110100000010101100000";
                        f_reg(317) <= "00010101100110101111111111111100";
                        f_reg(318) <= "10001100000111010000010110101100";
                        f_reg(319) <= "10001111101011010000010101100100";
                        f_reg(320) <= "10001100000111010000010110101100";
                        f_reg(321) <= "10001111101110110000010101100100";
                        f_reg(322) <= "00010101101110111111111111111100";
                        f_reg(323) <= "10001100000111010000010110101100";
                        f_reg(324) <= "10001111101011100000010101101000";
                        f_reg(325) <= "10001100000111010000010110101100";
                        f_reg(326) <= "10001111101111000000010101101000";
                        f_reg(327) <= "00010101110111001111111111111100";
                        f_reg(328) <= "10001100000111010000010110101100";
                        f_reg(329) <= "10001111101111100000010101101100";
                        f_reg(330) <= "10001100000111010000010110101100";
                        f_reg(331) <= "10001111101111110000010101101100";
                        f_reg(332) <= "00010111110111111111111111111100";
                        f_reg(333) <= "00010000000000001111111100111110";
                        f_reg(334) <= "00000000000000000000000000000000";
                        f_reg(335) <= "00000000000000000000000000000000";
                        f_reg(336) <= "00000000000000000000000000000000";
                        f_reg(337) <= "00000000000000000000000000000000";
                        f_reg(338) <= "00000000000000000000000000000000";
                        f_reg(339) <= "00000000000000000000000000000000";
                        f_reg(340) <= "00000000000000000000000000000000";
                        f_reg(341) <= "00000000000000000000000000000000";
                        f_reg(342) <= "00000000000000000000000000000000";
                        f_reg(343) <= "00000000000000000000000000000000";
                        f_reg(344) <= "00000000000000000000000000000000";
                        f_reg(345) <= "00000000000000000000000000000000";
                        f_reg(346) <= "00000000000000000000000000000000";
                        f_reg(347) <= "00000000000000000000000000000000";
                        f_reg(348) <= "00000000000000000000000000000000";
                        f_reg(349) <= "00000000000000000000000000000000";
                        f_reg(350) <= "00000000000000000000000000000000";
                        f_reg(351) <= "00000000000000000000000000000000";
                        f_reg(352) <= "00000000000000000000000000000000";
                        f_reg(353) <= "00000000000000000000000000000000";
                        f_reg(354) <= "00000000000000000000000000000000";
                        f_reg(355) <= "00000000000000000000000000000000";
                        f_reg(356) <= "00000000000000000000000000000000";
                        f_reg(357) <= "00000000000000000000000000000000";
                        f_reg(358) <= "00000000000000000000000000000000";
                        f_reg(359) <= "00000000000000000000000000000000";
                        f_reg(360) <= "00000000000000000000000000000000";
                        f_reg(361) <= "00000000000000000000000000000000";
                        f_reg(362) <= "00000000000000000000000000000000";
                        f_reg(363) <= "00000000000000000000000000000000";
                        f_reg(364) <= "00000000000000000000001111100111";
                        f_reg(365) <= "00000000000000000000000000000000";
                        f_reg(366) <= "00000000000000000000000000000000";
                        f_reg(367) <= "00000000000000000000000000000000";
                        f_reg(368) <= "00000000000000000000000000000000";
                        f_reg(369) <= "00000000000000000000000000000000";
                        f_reg(370) <= "00000000000000000000000000000000";
                        f_reg(371) <= "00000000000000000000000000000000";
                        f_reg(372) <= "00000000000000000000000000000000";
                        f_reg(373) <= "00000000000000000000000000000000";
                        f_reg(374) <= "00000000000000000000000000000000";
                        f_reg(375) <= "00000000000000000000000000000000";
                        f_reg(376) <= "00000000000000000000000000000000";
                        f_reg(377) <= "00000000000000000000000000000000";
                        f_reg(378) <= "00000000000000000000000000000000";
                        f_reg(379) <= "00000000000000000000000000000000";
                        f_reg(380) <= "00000000000000000000000000000000";
                        f_reg(381) <= "00000000000000000000000000000000";
                        f_reg(382) <= "00000000000000000000000000000000";
                        f_reg(383) <= "00000000000000000000000000000000";
                        f_reg(384) <= "00000000000000000000000000000000";
                        f_reg(385) <= "00000000000000000000000000000000";
                        f_reg(386) <= "00000000000000000000000000000000";
                        f_reg(387) <= "00000000000000000000000000000000";
                        f_reg(388) <= "00000000000000000000000000000000";
                        f_reg(389) <= "00000000000000000000000000000000";
                        f_reg(390) <= "00000000000000000000000000000000";
                        f_reg(391) <= "00000000000000000000000000000000";
                        f_reg(392) <= "00000000000000000000000000000000";
                        f_reg(393) <= "00000000000000000000000000000000";
                        f_reg(394) <= "00000000000000000000000000000000";
                        f_reg(395) <= "00000000000000000000000000000000";
                        f_reg(396) <= "00000000000000000000000000000000";
                        f_reg(397) <= "00000000000000000000000000000000";
                        f_reg(398) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011101010000101101";
                        f_reg(4) <= "00000000000000000001010011000011";
                        f_reg(5) <= "00000000000000100001110111000000";
                        f_reg(6) <= "00111000001001000010001100100111";
                        f_reg(7) <= "00000000001001000010100000100101";
                        f_reg(8) <= "00111000010001100000110100110100";
                        f_reg(9) <= "00101100011001110100011001001000";
                        f_reg(10) <= "00100100110010001111010001101010";
                        f_reg(11) <= "00000000110001010100100000000110";
                        f_reg(12) <= "00100001000010101000111000000001";
                        f_reg(13) <= "00000000000001010101100000000111";
                        f_reg(14) <= "00000000110001100110000000000100";
                        f_reg(15) <= "00110101001011010100110100111001";
                        f_reg(16) <= "00000000000011000111000010000011";
                        f_reg(17) <= "10101100000000100000001000111100";
                        f_reg(18) <= "00110001110011110111100111000111";
                        f_reg(19) <= "00000000000000000000000000000000";
                        f_reg(20) <= "00000000000000000000000000000000";
                        f_reg(21) <= "00101001001100001101011001101000";
                        f_reg(22) <= "10101100000001110000001001000000";
                        f_reg(23) <= "00000000000010111000110111000010";
                        f_reg(24) <= "00100110001100101011010101001001";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00111100000100111000101011001111";
                        f_reg(27) <= "00000000000000000000000000000000";
                        f_reg(28) <= "00000000000100111010010101000010";
                        f_reg(29) <= "00000001101101001010100000100011";
                        f_reg(30) <= "00110100011101100011000000000110";
                        f_reg(31) <= "10101100000010100000001001000100";
                        f_reg(32) <= "00100110000101111111011111011000";
                        f_reg(33) <= "00000000000101111100000110000011";
                        f_reg(34) <= "00000000000000000000000000000000";
                        f_reg(35) <= "10101100000101100000001001001000";
                        f_reg(36) <= "00000010101110001100100000100111";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "10101100000011110000001001001100";
                        f_reg(39) <= "00000010010110011101000000101011";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "10101100000100010000001001010000";
                        f_reg(42) <= "00000000000000000000000000000000";
                        f_reg(43) <= "10101100000110100000001001010100";
                        f_reg(44) <= "00100011111111111111111111111111";
                        f_reg(45) <= "00011111111000001111111111010110";
                        f_reg(46) <= "00010000000000000000000101100001";
                        f_reg(47) <= "00111100000111100000001111100111";
                        f_reg(48) <= "00111100000111110000001111100111";
                        f_reg(49) <= "00000000000111101111010000000010";
                        f_reg(50) <= "00000000000111111111110000000010";
                        f_reg(51) <= "00111100000000011101010000101101";
                        f_reg(52) <= "00111100000011111101010000101101";
                        f_reg(53) <= "00000000000000000001010011000011";
                        f_reg(54) <= "00000000000000001000010011000011";
                        f_reg(55) <= "00000000000000100001110111000000";
                        f_reg(56) <= "00000000000100001000110111000000";
                        f_reg(57) <= "00111000001001000010001100100111";
                        f_reg(58) <= "00111001111100100010001100100111";
                        f_reg(59) <= "00000000001001000010100000100101";
                        f_reg(60) <= "00000001111100101001100000100101";
                        f_reg(61) <= "00111000010001100000110100110100";
                        f_reg(62) <= "00111010000101000000110100110100";
                        f_reg(63) <= "00101100011001110100011001001000";
                        f_reg(64) <= "00101110001101010100011001001000";
                        f_reg(65) <= "00100100110010001111010001101010";
                        f_reg(66) <= "00100110100101101111010001101010";
                        f_reg(67) <= "00000000110001010100100000000110";
                        f_reg(68) <= "00000010100100111011100000000110";
                        f_reg(69) <= "00100001000010101000111000000001";
                        f_reg(70) <= "00100010110110001000111000000001";
                        f_reg(71) <= "00000000000001010101100000000111";
                        f_reg(72) <= "00000000000100111100100000000111";
                        f_reg(73) <= "00000000110001100110000000000100";
                        f_reg(74) <= "00000010100101001101000000000100";
                        f_reg(75) <= "00110101001011010100110100111001";
                        f_reg(76) <= "00110110111110110100110100111001";
                        f_reg(77) <= "00000000000011000111000010000011";
                        f_reg(78) <= "00000000000110101110000010000011";
                        f_reg(79) <= "00010100010100000000000010110011";
                        f_reg(80) <= "10101100000000100000001000111100";
                        f_reg(81) <= "00110001110000010111100111000111";
                        f_reg(82) <= "00110011100011110111100111000111";
                        f_reg(83) <= "00000000000000000000000000000000";
                        f_reg(84) <= "00000000000000000000000000000000";
                        f_reg(85) <= "00000000000000000000000000000000";
                        f_reg(86) <= "00000000000000000000000000000000";
                        f_reg(87) <= "00101001001001001101011001101000";
                        f_reg(88) <= "00101010111100101101011001101000";
                        f_reg(89) <= "00010100111101010000000010101001";
                        f_reg(90) <= "10101100000001110000001001000000";
                        f_reg(91) <= "00000000000010110100010111000010";
                        f_reg(92) <= "00000000000110011011010111000010";
                        f_reg(93) <= "00100101000001011011010101001001";
                        f_reg(94) <= "00100110110100111011010101001001";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000000000000000000000000000";
                        f_reg(97) <= "00111100000001101000101011001111";
                        f_reg(98) <= "00111100000101001000101011001111";
                        f_reg(99) <= "00000000000000000000000000000000";
                        f_reg(100) <= "00000000000000000000000000000000";
                        f_reg(101) <= "00000000000001100110010101000010";
                        f_reg(102) <= "00000000000101001101010101000010";
                        f_reg(103) <= "00000001101011000001000000100011";
                        f_reg(104) <= "00000011011110101000000000100011";
                        f_reg(105) <= "00110100011011100011000000000110";
                        f_reg(106) <= "00110110001111000011000000000110";
                        f_reg(107) <= "00010101010110000000000010010111";
                        f_reg(108) <= "10101100000010100000001001000100";
                        f_reg(109) <= "00100100100010011111011111011000";
                        f_reg(110) <= "00100110010101111111011111011000";
                        f_reg(111) <= "00000000000010010011100110000011";
                        f_reg(112) <= "00000000000101111010100110000011";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00010101110111000000000010001111";
                        f_reg(116) <= "10101100000011100000001001001000";
                        f_reg(117) <= "00000000010001110101100000100111";
                        f_reg(118) <= "00000010000101011100100000100111";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000000000000000000000000000";
                        f_reg(121) <= "00010100001011110000000010001001";
                        f_reg(122) <= "10101100000000010000001001001100";
                        f_reg(123) <= "00000000101010110011000000101011";
                        f_reg(124) <= "00000010011110011010000000101011";
                        f_reg(125) <= "00000000000000000000000000000000";
                        f_reg(126) <= "00000000000000000000000000000000";
                        f_reg(127) <= "00010101000101100000000010000011";
                        f_reg(128) <= "10101100000010000000001001010000";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010100110101000000000001111111";
                        f_reg(132) <= "10101100000001100000001001010100";
                        f_reg(133) <= "00100011110111011111111100000110";
                        f_reg(134) <= "00010011101000000000000000010001";
                        f_reg(135) <= "00100011110111011111111000001100";
                        f_reg(136) <= "00010011101000000000000000001111";
                        f_reg(137) <= "00100011110111011111110100010010";
                        f_reg(138) <= "00010011101000000000000000001101";
                        f_reg(139) <= "00100011110111101111111111111111";
                        f_reg(140) <= "00100011111111111111111111111111";
                        f_reg(141) <= "00010111110111110000000001110101";
                        f_reg(142) <= "00011111111000001111111110100101";
                        f_reg(143) <= "00010000000000000000000100000000";
                        f_reg(144) <= "00000000000000000000000000000000";
                        f_reg(145) <= "00000000000000000000000000000000";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000000000000000000000000000";
                        f_reg(149) <= "00000000000000000000000000000000";
                        f_reg(150) <= "00000000000000000000000000000000";
                        f_reg(151) <= "10001100000111010000010110101100";
                        f_reg(152) <= "00011111101000000000000000000011";
                        f_reg(153) <= "00100000000111010000000000111100";
                        f_reg(154) <= "00010000000000000000000000000010";
                        f_reg(155) <= "00100000000111010000000000000000";
                        f_reg(156) <= "00010100001011110000000001100110";
                        f_reg(157) <= "10101111101000010000010100110100";
                        f_reg(158) <= "10001100000111010000010110101100";
                        f_reg(159) <= "00011111101000000000000000000011";
                        f_reg(160) <= "00100000000111010000000000111100";
                        f_reg(161) <= "00010000000000000000000000000010";
                        f_reg(162) <= "00100000000111010000000000000000";
                        f_reg(163) <= "00010100010100000000000001011111";
                        f_reg(164) <= "10101111101000100000010100111000";
                        f_reg(165) <= "10001100000111010000010110101100";
                        f_reg(166) <= "00011111101000000000000000000011";
                        f_reg(167) <= "00100000000111010000000000111100";
                        f_reg(168) <= "00010000000000000000000000000010";
                        f_reg(169) <= "00100000000111010000000000000000";
                        f_reg(170) <= "00010100011100010000000001011000";
                        f_reg(171) <= "10101111101000110000010100111100";
                        f_reg(172) <= "10001100000111010000010110101100";
                        f_reg(173) <= "00011111101000000000000000000011";
                        f_reg(174) <= "00100000000111010000000000111100";
                        f_reg(175) <= "00010000000000000000000000000010";
                        f_reg(176) <= "00100000000111010000000000000000";
                        f_reg(177) <= "00010100100100100000000001010001";
                        f_reg(178) <= "10101111101001000000010101000000";
                        f_reg(179) <= "10001100000111010000010110101100";
                        f_reg(180) <= "00011111101000000000000000000011";
                        f_reg(181) <= "00100000000111010000000000111100";
                        f_reg(182) <= "00010000000000000000000000000010";
                        f_reg(183) <= "00100000000111010000000000000000";
                        f_reg(184) <= "00010100101100110000000001001010";
                        f_reg(185) <= "10101111101001010000010101000100";
                        f_reg(186) <= "10001100000111010000010110101100";
                        f_reg(187) <= "00011111101000000000000000000011";
                        f_reg(188) <= "00100000000111010000000000111100";
                        f_reg(189) <= "00010000000000000000000000000010";
                        f_reg(190) <= "00100000000111010000000000000000";
                        f_reg(191) <= "00010100110101000000000001000011";
                        f_reg(192) <= "10101111101001100000010101001000";
                        f_reg(193) <= "10001100000111010000010110101100";
                        f_reg(194) <= "00011111101000000000000000000011";
                        f_reg(195) <= "00100000000111010000000000111100";
                        f_reg(196) <= "00010000000000000000000000000010";
                        f_reg(197) <= "00100000000111010000000000000000";
                        f_reg(198) <= "00010100111101010000000000111100";
                        f_reg(199) <= "10101111101001110000010101001100";
                        f_reg(200) <= "10001100000111010000010110101100";
                        f_reg(201) <= "00011111101000000000000000000011";
                        f_reg(202) <= "00100000000111010000000000111100";
                        f_reg(203) <= "00010000000000000000000000000010";
                        f_reg(204) <= "00100000000111010000000000000000";
                        f_reg(205) <= "00010101000101100000000000110101";
                        f_reg(206) <= "10101111101010000000010101010000";
                        f_reg(207) <= "10001100000111010000010110101100";
                        f_reg(208) <= "00011111101000000000000000000011";
                        f_reg(209) <= "00100000000111010000000000111100";
                        f_reg(210) <= "00010000000000000000000000000010";
                        f_reg(211) <= "00100000000111010000000000000000";
                        f_reg(212) <= "00010101001101110000000000101110";
                        f_reg(213) <= "10101111101010010000010101010100";
                        f_reg(214) <= "10001100000111010000010110101100";
                        f_reg(215) <= "00011111101000000000000000000011";
                        f_reg(216) <= "00100000000111010000000000111100";
                        f_reg(217) <= "00010000000000000000000000000010";
                        f_reg(218) <= "00100000000111010000000000000000";
                        f_reg(219) <= "00010101010110000000000000100111";
                        f_reg(220) <= "10101111101010100000010101011000";
                        f_reg(221) <= "10001100000111010000010110101100";
                        f_reg(222) <= "00011111101000000000000000000011";
                        f_reg(223) <= "00100000000111010000000000111100";
                        f_reg(224) <= "00010000000000000000000000000010";
                        f_reg(225) <= "00100000000111010000000000000000";
                        f_reg(226) <= "00010101011110010000000000100000";
                        f_reg(227) <= "10101111101010110000010101011100";
                        f_reg(228) <= "10001100000111010000010110101100";
                        f_reg(229) <= "00011111101000000000000000000011";
                        f_reg(230) <= "00100000000111010000000000111100";
                        f_reg(231) <= "00010000000000000000000000000010";
                        f_reg(232) <= "00100000000111010000000000000000";
                        f_reg(233) <= "00010101100110100000000000011001";
                        f_reg(234) <= "10101111101011000000010101100000";
                        f_reg(235) <= "10001100000111010000010110101100";
                        f_reg(236) <= "00011111101000000000000000000011";
                        f_reg(237) <= "00100000000111010000000000111100";
                        f_reg(238) <= "00010000000000000000000000000010";
                        f_reg(239) <= "00100000000111010000000000000000";
                        f_reg(240) <= "00010101101110110000000000010010";
                        f_reg(241) <= "10101111101011010000010101100100";
                        f_reg(242) <= "10001100000111010000010110101100";
                        f_reg(243) <= "00011111101000000000000000000011";
                        f_reg(244) <= "00100000000111010000000000111100";
                        f_reg(245) <= "00010000000000000000000000000010";
                        f_reg(246) <= "00100000000111010000000000000000";
                        f_reg(247) <= "00010101110111000000000000001011";
                        f_reg(248) <= "10101111101011100000010101101000";
                        f_reg(249) <= "10001100000111010000010110101100";
                        f_reg(250) <= "00011111101000000000000000000011";
                        f_reg(251) <= "00100000000111010000000000111100";
                        f_reg(252) <= "00010000000000000000000000000010";
                        f_reg(253) <= "00100000000111010000000000000000";
                        f_reg(254) <= "00010111110111110000000000000100";
                        f_reg(255) <= "10101111101111100000010101101100";
                        f_reg(256) <= "10101100000111010000010110101100";
                        f_reg(257) <= "00010000000000001111111110001010";
                        f_reg(258) <= "10001100000111010000010110101100";
                        f_reg(259) <= "10001111101000010000010100110100";
                        f_reg(260) <= "10001100000111010000010110101100";
                        f_reg(261) <= "10001111101011110000010100110100";
                        f_reg(262) <= "00010100001011111111111111111100";
                        f_reg(263) <= "10001100000111010000010110101100";
                        f_reg(264) <= "10001111101000100000010100111000";
                        f_reg(265) <= "10001100000111010000010110101100";
                        f_reg(266) <= "10001111101100000000010100111000";
                        f_reg(267) <= "00010100010100001111111111111100";
                        f_reg(268) <= "10001100000111010000010110101100";
                        f_reg(269) <= "10001111101000110000010100111100";
                        f_reg(270) <= "10001100000111010000010110101100";
                        f_reg(271) <= "10001111101100010000010100111100";
                        f_reg(272) <= "00010100011100011111111111111100";
                        f_reg(273) <= "10001100000111010000010110101100";
                        f_reg(274) <= "10001111101001000000010101000000";
                        f_reg(275) <= "10001100000111010000010110101100";
                        f_reg(276) <= "10001111101100100000010101000000";
                        f_reg(277) <= "00010100100100101111111111111100";
                        f_reg(278) <= "10001100000111010000010110101100";
                        f_reg(279) <= "10001111101001010000010101000100";
                        f_reg(280) <= "10001100000111010000010110101100";
                        f_reg(281) <= "10001111101100110000010101000100";
                        f_reg(282) <= "00010100101100111111111111111100";
                        f_reg(283) <= "10001100000111010000010110101100";
                        f_reg(284) <= "10001111101001100000010101001000";
                        f_reg(285) <= "10001100000111010000010110101100";
                        f_reg(286) <= "10001111101101000000010101001000";
                        f_reg(287) <= "00010100110101001111111111111100";
                        f_reg(288) <= "10001100000111010000010110101100";
                        f_reg(289) <= "10001111101001110000010101001100";
                        f_reg(290) <= "10001100000111010000010110101100";
                        f_reg(291) <= "10001111101101010000010101001100";
                        f_reg(292) <= "00010100111101011111111111111100";
                        f_reg(293) <= "10001100000111010000010110101100";
                        f_reg(294) <= "10001111101010000000010101010000";
                        f_reg(295) <= "10001100000111010000010110101100";
                        f_reg(296) <= "10001111101101100000010101010000";
                        f_reg(297) <= "00010101000101101111111111111100";
                        f_reg(298) <= "10001100000111010000010110101100";
                        f_reg(299) <= "10001111101010010000010101010100";
                        f_reg(300) <= "10001100000111010000010110101100";
                        f_reg(301) <= "10001111101101110000010101010100";
                        f_reg(302) <= "00010101001101111111111111111100";
                        f_reg(303) <= "10001100000111010000010110101100";
                        f_reg(304) <= "10001111101010100000010101011000";
                        f_reg(305) <= "10001100000111010000010110101100";
                        f_reg(306) <= "10001111101110000000010101011000";
                        f_reg(307) <= "00010101010110001111111111111100";
                        f_reg(308) <= "10001100000111010000010110101100";
                        f_reg(309) <= "10001111101010110000010101011100";
                        f_reg(310) <= "10001100000111010000010110101100";
                        f_reg(311) <= "10001111101110010000010101011100";
                        f_reg(312) <= "00010101011110011111111111111100";
                        f_reg(313) <= "10001100000111010000010110101100";
                        f_reg(314) <= "10001111101011000000010101100000";
                        f_reg(315) <= "10001100000111010000010110101100";
                        f_reg(316) <= "10001111101110100000010101100000";
                        f_reg(317) <= "00010101100110101111111111111100";
                        f_reg(318) <= "10001100000111010000010110101100";
                        f_reg(319) <= "10001111101011010000010101100100";
                        f_reg(320) <= "10001100000111010000010110101100";
                        f_reg(321) <= "10001111101110110000010101100100";
                        f_reg(322) <= "00010101101110111111111111111100";
                        f_reg(323) <= "10001100000111010000010110101100";
                        f_reg(324) <= "10001111101011100000010101101000";
                        f_reg(325) <= "10001100000111010000010110101100";
                        f_reg(326) <= "10001111101111000000010101101000";
                        f_reg(327) <= "00010101110111001111111111111100";
                        f_reg(328) <= "10001100000111010000010110101100";
                        f_reg(329) <= "10001111101111100000010101101100";
                        f_reg(330) <= "10001100000111010000010110101100";
                        f_reg(331) <= "10001111101111110000010101101100";
                        f_reg(332) <= "00010111110111111111111111111100";
                        f_reg(333) <= "00010000000000001111111100111110";
                        f_reg(334) <= "00000000000000000000000000000000";
                        f_reg(335) <= "00000000000000000000000000000000";
                        f_reg(336) <= "00000000000000000000000000000000";
                        f_reg(337) <= "00000000000000000000000000000000";
                        f_reg(338) <= "00000000000000000000000000000000";
                        f_reg(339) <= "00000000000000000000000000000000";
                        f_reg(340) <= "00000000000000000000000000000000";
                        f_reg(341) <= "00000000000000000000000000000000";
                        f_reg(342) <= "00000000000000000000000000000000";
                        f_reg(343) <= "00000000000000000000000000000000";
                        f_reg(344) <= "00000000000000000000000000000000";
                        f_reg(345) <= "00000000000000000000000000000000";
                        f_reg(346) <= "00000000000000000000000000000000";
                        f_reg(347) <= "00000000000000000000000000000000";
                        f_reg(348) <= "00000000000000000000000000000000";
                        f_reg(349) <= "00000000000000000000000000000000";
                        f_reg(350) <= "00000000000000000000000000000000";
                        f_reg(351) <= "00000000000000000000000000000000";
                        f_reg(352) <= "00000000000000000000000000000000";
                        f_reg(353) <= "00000000000000000000000000000000";
                        f_reg(354) <= "00000000000000000000000000000000";
                        f_reg(355) <= "00000000000000000000000000000000";
                        f_reg(356) <= "00000000000000000000000000000000";
                        f_reg(357) <= "00000000000000000000000000000000";
                        f_reg(358) <= "00000000000000000000000000000000";
                        f_reg(359) <= "00000000000000000000000000000000";
                        f_reg(360) <= "00000000000000000000000000000000";
                        f_reg(361) <= "00000000000000000000000000000000";
                        f_reg(362) <= "00000000000000000000000000000000";
                        f_reg(363) <= "00000000000000000000000000000000";
                        f_reg(364) <= "00000000000000000000001111100111";
                        f_reg(365) <= "00000000000000000000000000000000";
                        f_reg(366) <= "00000000000000000000000000000000";
                        f_reg(367) <= "00000000000000000000000000000000";
                        f_reg(368) <= "00000000000000000000000000000000";
                        f_reg(369) <= "00000000000000000000000000000000";
                        f_reg(370) <= "00000000000000000000000000000000";
                        f_reg(371) <= "00000000000000000000000000000000";
                        f_reg(372) <= "00000000000000000000000000000000";
                        f_reg(373) <= "00000000000000000000000000000000";
                        f_reg(374) <= "00000000000000000000000000000000";
                        f_reg(375) <= "00000000000000000000000000000000";
                        f_reg(376) <= "00000000000000000000000000000000";
                        f_reg(377) <= "00000000000000000000000000000000";
                        f_reg(378) <= "00000000000000000000000000000000";
                        f_reg(379) <= "00000000000000000000000000000000";
                        f_reg(380) <= "00000000000000000000000000000000";
                        f_reg(381) <= "00000000000000000000000000000000";
                        f_reg(382) <= "00000000000000000000000000000000";
                        f_reg(383) <= "00000000000000000000000000000000";
                        f_reg(384) <= "00000000000000000000000000000000";
                        f_reg(385) <= "00000000000000000000000000000000";
                        f_reg(386) <= "00000000000000000000000000000000";
                        f_reg(387) <= "00000000000000000000000000000000";
                        f_reg(388) <= "00000000000000000000000000000000";
                        f_reg(389) <= "00000000000000000000000000000000";
                        f_reg(390) <= "00000000000000000000000000000000";
                        f_reg(391) <= "00000000000000000000000000000000";
                        f_reg(392) <= "00000000000000000000000000000000";
                        f_reg(393) <= "00000000000000000000000000000000";
                        f_reg(394) <= "00000000000000000000000000000000";
                        f_reg(395) <= "00000000000000000000000000000000";
                        f_reg(396) <= "00000000000000000000000000000000";
                        f_reg(397) <= "00000000000000000000000000000000";
                        f_reg(398) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test31_Reg_COMBINED;
