--| Test73_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:13:08
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test73_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test73_Reg_COMBINED;

architecture a_Test73_Reg_COMBINED of Test73_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 496) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 496) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100");--  495 - 1980

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000010011010011001001", --    2 -    8
      "00111100000000101001011011000110", --    3 -   12
      "00000000000000010001100000000110", --    4 -   16
      "00101000001001000101110010010011", --    5 -   20
      "10101100000001000000001110101000", --    6 -   24
      "00000000000000000010100000100100", --    7 -   28
      "00000000001000000011000000000110", --    8 -   32
      "00000000110000010011100000100101", --    9 -   36
      "00000000000000000000000000000000", --   10 -   40
      "00000000110000000100000000100010", --   11 -   44
      "00000000000010000100110101000000", --   12 -   48
      "00100100101010101101000010011100", --   13 -   52
      "00000001010001010101100000100011", --   14 -   56
      "00101001011011000011010101010101", --   15 -   60
      "00000000011001000110100000100110", --   16 -   64
      "00000001100001100111000000101010", --   17 -   68
      "00101001110011111011100100100011", --   18 -   72
      "00000000001010111000000000000111", --   19 -   76
      "10101100000010000000001110101100", --   20 -   80
      "00000001101001111000100000000100", --   21 -   84
      "00000000000000000000000000000000", --   22 -   88
      "00000000010000011001000000100101", --   23 -   92
      "00000001011011001001100000100010", --   24 -   96
      "10101100000000100000001110110000", --   25 -  100
      "00000001100011011010000000100101", --   26 -  104
      "00000000000100111010111101000010", --   27 -  108
      "00000010010001111011000000100100", --   28 -  112
      "00110001001101110111010101110011", --   29 -  116
      "00000000000011101100011011000011", --   30 -  120
      "00000000010101011100100000000110", --   31 -  124
      "00000010100001011101000000100011", --   32 -  128
      "00111001110110111101011111110100", --   33 -  132
      "00000000000000000000000000000000", --   34 -  136
      "00000000010100101110000000101010", --   35 -  140
      "10101100000110100000001110110100", --   36 -  144
      "00000010101101101110100000100000", --   37 -  148
      "00000010001010001111000000100110", --   38 -  152
      "00000010000110010101000000100101", --   39 -  156
      "00000011100110000001100000100001", --   40 -  160
      "00000000011010100010000000100000", --   41 -  164
      "00000000000101000011001110000000", --   42 -  168
      "00000010110110000000100000100100", --   43 -  172
      "00000001111111010101100000100110", --   44 -  176
      "00000000000000000000000000000000", --   45 -  180
      "00111100000011011000001101011100", --   46 -  184
      "00000010111110011001100000100100", --   47 -  188
      "00000001010110000011100000100010", --   48 -  192
      "00000001100001100100100000000111", --   49 -  196
      "00000001001001000010100000100011", --   50 -  200
      "10101100000110110000001110111000", --   51 -  204
      "00000000111100110111000000100101", --   52 -  208
      "10101100000011100000001110111100", --   53 -  212
      "00000000000001010001000001000000", --   54 -  216
      "00110011110100101010011101011010", --   55 -  220
      "00000001011000101101000000000111", --   56 -  224
      "00000000000000011010110111000000", --   57 -  228
      "00000011101110001000100000101011", --   58 -  232
      "00000010101110100100000000000110", --   59 -  236
      "00100101101100000110000001101101", --   60 -  240
      "00000000000000000000000000000000", --   61 -  244
      "00000000000000000000000000000000", --   62 -  248
      "00000000000000000000000000000000", --   63 -  252
      "00000000000000000000000000000000", --   64 -  256
      "10101100000100000000001111000000", --   65 -  260
      "10101100000100010000001111000100", --   66 -  264
      "10101100000111010000001111001000", --   67 -  268
      "10101100000010000000001111001100", --   68 -  272
      "10101100000100100000001111010000", --   69 -  276
      "00100011111111111111111111111111", --   70 -  280
      "00011111111000001111111110111011", --   71 -  284
      "00010000000000000000000110100111", --   72 -  288
      "00111100000111100000001111100111", --   73 -  292
      "00111100000111110000001111100111", --   74 -  296
      "00000000000111101111010000000010", --   75 -  300
      "00000000000111111111110000000010", --   76 -  304
      "00111100000000010011010011001001", --   77 -  308
      "00111100000011110011010011001001", --   78 -  312
      "00111100000000101001011011000110", --   79 -  316
      "00111100000100001001011011000110", --   80 -  320
      "00000000000000010001100000000110", --   81 -  324
      "00000000000011111000100000000110", --   82 -  328
      "00101000001001000101110010010011", --   83 -  332
      "00101001111100100101110010010011", --   84 -  336
      "00010100100100100000000100001101", --   85 -  340
      "10101100000001000000001110101000", --   86 -  344
      "00000000000000000010100000100100", --   87 -  348
      "00000000000000001001100000100100", --   88 -  352
      "00000000001000000011000000000110", --   89 -  356
      "00000001111000001010000000000110", --   90 -  360
      "00000000110000010011100000100101", --   91 -  364
      "00000010100011111010100000100101", --   92 -  368
      "00000000000000000000000000000000", --   93 -  372
      "00000000000000000000000000000000", --   94 -  376
      "00000000110000000100000000100010", --   95 -  380
      "00000010100000001011000000100010", --   96 -  384
      "00000000000010000100110101000000", --   97 -  388
      "00000000000101101011110101000000", --   98 -  392
      "00100100101010101101000010011100", --   99 -  396
      "00100110011110001101000010011100", --  100 -  400
      "00000001010001010101100000100011", --  101 -  404
      "00000011000100111100100000100011", --  102 -  408
      "00101001011011000011010101010101", --  103 -  412
      "00101011001110100011010101010101", --  104 -  416
      "00000000011001000110100000100110", --  105 -  420
      "00000010001100101101100000100110", --  106 -  424
      "00000001100001100111000000101010", --  107 -  428
      "00000011010101001110000000101010", --  108 -  432
      "00101001110010101011100100100011", --  109 -  436
      "00101011100110001011100100100011", --  110 -  440
      "00000000001010110001100000000111", --  111 -  444
      "00000001111110011000100000000111", --  112 -  448
      "00010101000101100000000011110001", --  113 -  452
      "10101100000010000000001110101100", --  114 -  456
      "00000001101001110010000000000100", --  115 -  460
      "00000011011101011001000000000100", --  116 -  464
      "00000000000000000000000000000000", --  117 -  468
      "00000000000000000000000000000000", --  118 -  472
      "00000000010000010011000000100101", --  119 -  476
      "00000010000011111010000000100101", --  120 -  480
      "00000001011011000000100000100010", --  121 -  484
      "00000011001110100111100000100010", --  122 -  488
      "00010100010100000000000011100111", --  123 -  492
      "10101100000000100000001110110000", --  124 -  496
      "00000001100011010101100000100101", --  125 -  500
      "00000011010110111100100000100101", --  126 -  504
      "00000000000000010110111101000010", --  127 -  508
      "00000000000011111101111101000010", --  128 -  512
      "00000000110001110000100000100100", --  129 -  516
      "00000010100101010111100000100100", --  130 -  520
      "00110001001001110111010101110011", --  131 -  524
      "00110010111101010111010101110011", --  132 -  528
      "00000000000011100100111011000011", --  133 -  532
      "00000000000111001011111011000011", --  134 -  536
      "00010101001101110000000011011011", --  135 -  540
      "10101100000010010000001111010100", --  136 -  544
      "00000000010011010100100000000110", --  137 -  548
      "00000010000110111011100000000110", --  138 -  552
      "00010101100110100000000011010111", --  139 -  556
      "10101100000011000000001111011000", --  140 -  560
      "00000001011001010110000000100011", --  141 -  564
      "00000011001100111101000000100011", --  142 -  568
      "00111001110001011101011111110100", --  143 -  572
      "00111011100100111101011111110100", --  144 -  576
      "00000000000000000000000000000000", --  145 -  580
      "00000000000000000000000000000000", --  146 -  584
      "00000000010001100111000000101010", --  147 -  588
      "00000010000101001110000000101010", --  148 -  592
      "00010101100110100000000011001101", --  149 -  596
      "10101100000011000000001110110100", --  150 -  600
      "00000001101000010001000000100000", --  151 -  604
      "00000011011011111000000000100000", --  152 -  608
      "00000000100010000011000000100110", --  153 -  612
      "00000010010101101010000000100110", --  154 -  616
      "00000000011010010110000000100101", --  155 -  620
      "00000010001101111101000000100101", --  156 -  624
      "10001100000011010000001111010100", --  157 -  628
      "10001100000110110000001111010100", --  158 -  632
      "00010101101110111111111111111110", --  159 -  636
      "00000001110011010010000000100001", --  160 -  640
      "00000011100110111001000000100001", --  161 -  644
      "00000000100011000100000000100000", --  162 -  648
      "00000010010110101011000000100000", --  163 -  652
      "00000000000010110001101110000000", --  164 -  656
      "00000000000110011000101110000000", --  165 -  660
      "00000000001011010111000000100100", --  166 -  664
      "00000001111110111110000000100100", --  167 -  668
      "00000001010000100010000000100110", --  168 -  672
      "00000011000100001001000000100110", --  169 -  676
      "00000000000000000000000000000000", --  170 -  680
      "00000000000000000000000000000000", --  171 -  684
      "00111100000010111000001101011100", --  172 -  688
      "00111100000110011000001101011100", --  173 -  692
      "00000000111010010000100000100100", --  174 -  696
      "00000010101101110111100000100100", --  175 -  700
      "00000001100011010101000000100010", --  176 -  704
      "00000011010110111100000000100010", --  177 -  708
      "10001100000001110000001111011000", --  178 -  712
      "10001100000101010000001111011000", --  179 -  716
      "00010100111101011111111111111110", --  180 -  720
      "00000000111000110100100000000111", --  181 -  724
      "00000010101100011011100000000111", --  182 -  728
      "00000001001010000110000000100011", --  183 -  732
      "00000010111101101101000000100011", --  184 -  736
      "00010100101100110000000010101001", --  185 -  740
      "10101100000001010000001110111000", --  186 -  744
      "00000001010000010001100000100101", --  187 -  748
      "00000011000011111000100000100101", --  188 -  752
      "00010100011100010000000010100101", --  189 -  756
      "10101100000000110000001110111100", --  190 -  760
      "00000000000011000011100001000000", --  191 -  764
      "00000000000110101010100001000000", --  192 -  768
      "00110000110010011010011101011010", --  193 -  772
      "00110010100101111010011101011010", --  194 -  776
      "00000000100001110100000000000111", --  195 -  780
      "00000010010101011011000000000111", --  196 -  784
      "00000000000011100010110111000000", --  197 -  788
      "00000000000111001001110111000000", --  198 -  792
      "00000000010011010101000000101011", --  199 -  796
      "00000010000110111100000000101011", --  200 -  800
      "00000000101010000000100000000110", --  201 -  804
      "00000010011101100111100000000110", --  202 -  808
      "00100101011000110110000001101101", --  203 -  812
      "00100111001100010110000001101101", --  204 -  816
      "00000000000000000000000000000000", --  205 -  820
      "00000000000000000000000000000000", --  206 -  824
      "00000000000000000000000000000000", --  207 -  828
      "00000000000000000000000000000000", --  208 -  832
      "00000000000000000000000000000000", --  209 -  836
      "00000000000000000000000000000000", --  210 -  840
      "00000000000000000000000000000000", --  211 -  844
      "00000000000000000000000000000000", --  212 -  848
      "00010100011100010000000010001101", --  213 -  852
      "10101100000000110000001111000000", --  214 -  856
      "00010101010110000000000010001011", --  215 -  860
      "10101100000010100000001111000100", --  216 -  864
      "00010100010100000000000010001001", --  217 -  868
      "10101100000000100000001111001000", --  218 -  872
      "00010100001011110000000010000111", --  219 -  876
      "10101100000000010000001111001100", --  220 -  880
      "00010101001101110000000010000101", --  221 -  884
      "10101100000010010000001111010000", --  222 -  888
      "00100011110111011111111100000110", --  223 -  892
      "00010011101000000000000000010111", --  224 -  896
      "00100011110111011111111000001100", --  225 -  900
      "00010011101000000000000000010101", --  226 -  904
      "00100011110111011111110100010010", --  227 -  908
      "00010011101000000000000000010011", --  228 -  912
      "00100011110111101111111111111111", --  229 -  916
      "00100011111111111111111111111111", --  230 -  920
      "00010111110111110000000001111011", --  231 -  924
      "00011111111000001111111101100101", --  232 -  928
      "00010000000000000000000100000110", --  233 -  932
      "00000000000000000000000000000000", --  234 -  936
      "00000000000000000000000000000000", --  235 -  940
      "00000000000000000000000000000000", --  236 -  944
      "00000000000000000000000000000000", --  237 -  948
      "00000000000000000000000000000000", --  238 -  952
      "00000000000000000000000000000000", --  239 -  956
      "00000000000000000000000000000000", --  240 -  960
      "00000000000000000000000000000000", --  241 -  964
      "00000000000000000000000000000000", --  242 -  968
      "00000000000000000000000000000000", --  243 -  972
      "00000000000000000000000000000000", --  244 -  976
      "00000000000000000000000000000000", --  245 -  980
      "00000000000000000000000000000000", --  246 -  984
      "10001100000111010000011100110000", --  247 -  988
      "00011111101000000000000000000011", --  248 -  992
      "00100000000111010000000000111100", --  249 -  996
      "00010000000000000000000000000010", --  250 - 1000
      "00100000000111010000000000000000", --  251 - 1004
      "00010100001011110000000001100110", --  252 - 1008
      "10101111101000010000011010111000", --  253 - 1012
      "10001100000111010000011100110000", --  254 - 1016
      "00011111101000000000000000000011", --  255 - 1020
      "00100000000111010000000000111100", --  256 - 1024
      "00010000000000000000000000000010", --  257 - 1028
      "00100000000111010000000000000000", --  258 - 1032
      "00010100010100000000000001011111", --  259 - 1036
      "10101111101000100000011010111100", --  260 - 1040
      "10001100000111010000011100110000", --  261 - 1044
      "00011111101000000000000000000011", --  262 - 1048
      "00100000000111010000000000111100", --  263 - 1052
      "00010000000000000000000000000010", --  264 - 1056
      "00100000000111010000000000000000", --  265 - 1060
      "00010100011100010000000001011000", --  266 - 1064
      "10101111101000110000011011000000", --  267 - 1068
      "10001100000111010000011100110000", --  268 - 1072
      "00011111101000000000000000000011", --  269 - 1076
      "00100000000111010000000000111100", --  270 - 1080
      "00010000000000000000000000000010", --  271 - 1084
      "00100000000111010000000000000000", --  272 - 1088
      "00010100100100100000000001010001", --  273 - 1092
      "10101111101001000000011011000100", --  274 - 1096
      "10001100000111010000011100110000", --  275 - 1100
      "00011111101000000000000000000011", --  276 - 1104
      "00100000000111010000000000111100", --  277 - 1108
      "00010000000000000000000000000010", --  278 - 1112
      "00100000000111010000000000000000", --  279 - 1116
      "00010100101100110000000001001010", --  280 - 1120
      "10101111101001010000011011001000", --  281 - 1124
      "10001100000111010000011100110000", --  282 - 1128
      "00011111101000000000000000000011", --  283 - 1132
      "00100000000111010000000000111100", --  284 - 1136
      "00010000000000000000000000000010", --  285 - 1140
      "00100000000111010000000000000000", --  286 - 1144
      "00010100110101000000000001000011", --  287 - 1148
      "10101111101001100000011011001100", --  288 - 1152
      "10001100000111010000011100110000", --  289 - 1156
      "00011111101000000000000000000011", --  290 - 1160
      "00100000000111010000000000111100", --  291 - 1164
      "00010000000000000000000000000010", --  292 - 1168
      "00100000000111010000000000000000", --  293 - 1172
      "00010100111101010000000000111100", --  294 - 1176
      "10101111101001110000011011010000", --  295 - 1180
      "10001100000111010000011100110000", --  296 - 1184
      "00011111101000000000000000000011", --  297 - 1188
      "00100000000111010000000000111100", --  298 - 1192
      "00010000000000000000000000000010", --  299 - 1196
      "00100000000111010000000000000000", --  300 - 1200
      "00010101000101100000000000110101", --  301 - 1204
      "10101111101010000000011011010100", --  302 - 1208
      "10001100000111010000011100110000", --  303 - 1212
      "00011111101000000000000000000011", --  304 - 1216
      "00100000000111010000000000111100", --  305 - 1220
      "00010000000000000000000000000010", --  306 - 1224
      "00100000000111010000000000000000", --  307 - 1228
      "00010101001101110000000000101110", --  308 - 1232
      "10101111101010010000011011011000", --  309 - 1236
      "10001100000111010000011100110000", --  310 - 1240
      "00011111101000000000000000000011", --  311 - 1244
      "00100000000111010000000000111100", --  312 - 1248
      "00010000000000000000000000000010", --  313 - 1252
      "00100000000111010000000000000000", --  314 - 1256
      "00010101010110000000000000100111", --  315 - 1260
      "10101111101010100000011011011100", --  316 - 1264
      "10001100000111010000011100110000", --  317 - 1268
      "00011111101000000000000000000011", --  318 - 1272
      "00100000000111010000000000111100", --  319 - 1276
      "00010000000000000000000000000010", --  320 - 1280
      "00100000000111010000000000000000", --  321 - 1284
      "00010101011110010000000000100000", --  322 - 1288
      "10101111101010110000011011100000", --  323 - 1292
      "10001100000111010000011100110000", --  324 - 1296
      "00011111101000000000000000000011", --  325 - 1300
      "00100000000111010000000000111100", --  326 - 1304
      "00010000000000000000000000000010", --  327 - 1308
      "00100000000111010000000000000000", --  328 - 1312
      "00010101100110100000000000011001", --  329 - 1316
      "10101111101011000000011011100100", --  330 - 1320
      "10001100000111010000011100110000", --  331 - 1324
      "00011111101000000000000000000011", --  332 - 1328
      "00100000000111010000000000111100", --  333 - 1332
      "00010000000000000000000000000010", --  334 - 1336
      "00100000000111010000000000000000", --  335 - 1340
      "00010101101110110000000000010010", --  336 - 1344
      "10101111101011010000011011101000", --  337 - 1348
      "10001100000111010000011100110000", --  338 - 1352
      "00011111101000000000000000000011", --  339 - 1356
      "00100000000111010000000000111100", --  340 - 1360
      "00010000000000000000000000000010", --  341 - 1364
      "00100000000111010000000000000000", --  342 - 1368
      "00010101110111000000000000001011", --  343 - 1372
      "10101111101011100000011011101100", --  344 - 1376
      "10001100000111010000011100110000", --  345 - 1380
      "00011111101000000000000000000011", --  346 - 1384
      "00100000000111010000000000111100", --  347 - 1388
      "00010000000000000000000000000010", --  348 - 1392
      "00100000000111010000000000000000", --  349 - 1396
      "00010111110111110000000000000100", --  350 - 1400
      "10101111101111100000011011110000", --  351 - 1404
      "10101100000111010000011100110000", --  352 - 1408
      "00010000000000001111111110000100", --  353 - 1412
      "10001100000111010000011100110000", --  354 - 1416
      "10001111101000010000011010111000", --  355 - 1420
      "10001100000111010000011100110000", --  356 - 1424
      "10001111101011110000011010111000", --  357 - 1428
      "00010100001011111111111111111100", --  358 - 1432
      "10001100000111010000011100110000", --  359 - 1436
      "10001111101000100000011010111100", --  360 - 1440
      "10001100000111010000011100110000", --  361 - 1444
      "10001111101100000000011010111100", --  362 - 1448
      "00010100010100001111111111111100", --  363 - 1452
      "10001100000111010000011100110000", --  364 - 1456
      "10001111101000110000011011000000", --  365 - 1460
      "10001100000111010000011100110000", --  366 - 1464
      "10001111101100010000011011000000", --  367 - 1468
      "00010100011100011111111111111100", --  368 - 1472
      "10001100000111010000011100110000", --  369 - 1476
      "10001111101001000000011011000100", --  370 - 1480
      "10001100000111010000011100110000", --  371 - 1484
      "10001111101100100000011011000100", --  372 - 1488
      "00010100100100101111111111111100", --  373 - 1492
      "10001100000111010000011100110000", --  374 - 1496
      "10001111101001010000011011001000", --  375 - 1500
      "10001100000111010000011100110000", --  376 - 1504
      "10001111101100110000011011001000", --  377 - 1508
      "00010100101100111111111111111100", --  378 - 1512
      "10001100000111010000011100110000", --  379 - 1516
      "10001111101001100000011011001100", --  380 - 1520
      "10001100000111010000011100110000", --  381 - 1524
      "10001111101101000000011011001100", --  382 - 1528
      "00010100110101001111111111111100", --  383 - 1532
      "10001100000111010000011100110000", --  384 - 1536
      "10001111101001110000011011010000", --  385 - 1540
      "10001100000111010000011100110000", --  386 - 1544
      "10001111101101010000011011010000", --  387 - 1548
      "00010100111101011111111111111100", --  388 - 1552
      "10001100000111010000011100110000", --  389 - 1556
      "10001111101010000000011011010100", --  390 - 1560
      "10001100000111010000011100110000", --  391 - 1564
      "10001111101101100000011011010100", --  392 - 1568
      "00010101000101101111111111111100", --  393 - 1572
      "10001100000111010000011100110000", --  394 - 1576
      "10001111101010010000011011011000", --  395 - 1580
      "10001100000111010000011100110000", --  396 - 1584
      "10001111101101110000011011011000", --  397 - 1588
      "00010101001101111111111111111100", --  398 - 1592
      "10001100000111010000011100110000", --  399 - 1596
      "10001111101010100000011011011100", --  400 - 1600
      "10001100000111010000011100110000", --  401 - 1604
      "10001111101110000000011011011100", --  402 - 1608
      "00010101010110001111111111111100", --  403 - 1612
      "10001100000111010000011100110000", --  404 - 1616
      "10001111101010110000011011100000", --  405 - 1620
      "10001100000111010000011100110000", --  406 - 1624
      "10001111101110010000011011100000", --  407 - 1628
      "00010101011110011111111111111100", --  408 - 1632
      "10001100000111010000011100110000", --  409 - 1636
      "10001111101011000000011011100100", --  410 - 1640
      "10001100000111010000011100110000", --  411 - 1644
      "10001111101110100000011011100100", --  412 - 1648
      "00010101100110101111111111111100", --  413 - 1652
      "10001100000111010000011100110000", --  414 - 1656
      "10001111101011010000011011101000", --  415 - 1660
      "10001100000111010000011100110000", --  416 - 1664
      "10001111101110110000011011101000", --  417 - 1668
      "00010101101110111111111111111100", --  418 - 1672
      "10001100000111010000011100110000", --  419 - 1676
      "10001111101011100000011011101100", --  420 - 1680
      "10001100000111010000011100110000", --  421 - 1684
      "10001111101111000000011011101100", --  422 - 1688
      "00010101110111001111111111111100", --  423 - 1692
      "10001100000111010000011100110000", --  424 - 1696
      "10001111101111100000011011110000", --  425 - 1700
      "10001100000111010000011100110000", --  426 - 1704
      "10001111101111110000011011110000", --  427 - 1708
      "00010111110111111111111111111100", --  428 - 1712
      "00010000000000001111111100111000", --  429 - 1716
      "00000000000000000000000000000000", --  430 - 1720
      "00000000000000000000000000000000", --  431 - 1724
      "00000000000000000000000000000000", --  432 - 1728
      "00000000000000000000000000000000", --  433 - 1732
      "00000000000000000000000000000000", --  434 - 1736
      "00000000000000000000000000000000", --  435 - 1740
      "00000000000000000000000000000000", --  436 - 1744
      "00000000000000000000000000000000", --  437 - 1748
      "00000000000000000000000000000000", --  438 - 1752
      "00000000000000000000000000000000", --  439 - 1756
      "00000000000000000000000000000000", --  440 - 1760
      "00000000000000000000000000000000", --  441 - 1764
      "00000000000000000000000000000000", --  442 - 1768
      "00000000000000000000000000000000", --  443 - 1772
      "00000000000000000000000000000000", --  444 - 1776
      "00000000000000000000000000000000", --  445 - 1780
      "00000000000000000000000000000000", --  446 - 1784
      "00000000000000000000000000000000", --  447 - 1788
      "00000000000000000000000000000000", --  448 - 1792
      "00000000000000000000000000000000", --  449 - 1796
      "00000000000000000000000000000000", --  450 - 1800
      "00000000000000000000000000000000", --  451 - 1804
      "00000000000000000000000000000000", --  452 - 1808
      "00000000000000000000000000000000", --  453 - 1812
      "00000000000000000000000000000000", --  454 - 1816
      "00000000000000000000000000000000", --  455 - 1820
      "00000000000000000000000000000000", --  456 - 1824
      "00000000000000000000000000000000", --  457 - 1828
      "00000000000000000000000000000000", --  458 - 1832
      "00000000000000000000000000000000", --  459 - 1836
      "00000000000000000000001111100111", --  460 - 1840
      "00000000000000000000000000000000", --  461 - 1844
      "00000000000000000000000000000000", --  462 - 1848
      "00000000000000000000000000000000", --  463 - 1852
      "00000000000000000000000000000000", --  464 - 1856
      "00000000000000000000000000000000", --  465 - 1860
      "00000000000000000000000000000000", --  466 - 1864
      "00000000000000000000000000000000", --  467 - 1868
      "00000000000000000000000000000000", --  468 - 1872
      "00000000000000000000000000000000", --  469 - 1876
      "00000000000000000000000000000000", --  470 - 1880
      "00000000000000000000000000000000", --  471 - 1884
      "00000000000000000000000000000000", --  472 - 1888
      "00000000000000000000000000000000", --  473 - 1892
      "00000000000000000000000000000000", --  474 - 1896
      "00000000000000000000000000000000", --  475 - 1900
      "00000000000000000000000000000000", --  476 - 1904
      "00000000000000000000000000000000", --  477 - 1908
      "00000000000000000000000000000000", --  478 - 1912
      "00000000000000000000000000000000", --  479 - 1916
      "00000000000000000000000000000000", --  480 - 1920
      "00000000000000000000000000000000", --  481 - 1924
      "00000000000000000000000000000000", --  482 - 1928
      "00000000000000000000000000000000", --  483 - 1932
      "00000000000000000000000000000000", --  484 - 1936
      "00000000000000000000000000000000", --  485 - 1940
      "00000000000000000000000000000000", --  486 - 1944
      "00000000000000000000000000000000", --  487 - 1948
      "00000000000000000000000000000000", --  488 - 1952
      "00000000000000000000000000000000", --  489 - 1956
      "00000000000000000000000000000000", --  490 - 1960
      "00000000000000000000000000000000", --  491 - 1964
      "00000000000000000000000000000000", --  492 - 1968
      "00000000000000000000000000000000", --  493 - 1972
      "00000000000000000000000000000000", --  494 - 1976
      "00000000000000000000000000000000");--  495 - 1980

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000010011010011001001";
         f_reg(4) <= "00111100000000101001011011000110";
         f_reg(5) <= "00000000000000010001100000000110";
         f_reg(6) <= "00101000001001000101110010010011";
         f_reg(7) <= "10101100000001000000001110101000";
         f_reg(8) <= "00000000000000000010100000100100";
         f_reg(9) <= "00000000001000000011000000000110";
         f_reg(10) <= "00000000110000010011100000100101";
         f_reg(11) <= "00000000000000000000000000000000";
         f_reg(12) <= "00000000110000000100000000100010";
         f_reg(13) <= "00000000000010000100110101000000";
         f_reg(14) <= "00100100101010101101000010011100";
         f_reg(15) <= "00000001010001010101100000100011";
         f_reg(16) <= "00101001011011000011010101010101";
         f_reg(17) <= "00000000011001000110100000100110";
         f_reg(18) <= "00000001100001100111000000101010";
         f_reg(19) <= "00101001110011111011100100100011";
         f_reg(20) <= "00000000001010111000000000000111";
         f_reg(21) <= "10101100000010000000001110101100";
         f_reg(22) <= "00000001101001111000100000000100";
         f_reg(23) <= "00000000000000000000000000000000";
         f_reg(24) <= "00000000010000011001000000100101";
         f_reg(25) <= "00000001011011001001100000100010";
         f_reg(26) <= "10101100000000100000001110110000";
         f_reg(27) <= "00000001100011011010000000100101";
         f_reg(28) <= "00000000000100111010111101000010";
         f_reg(29) <= "00000010010001111011000000100100";
         f_reg(30) <= "00110001001101110111010101110011";
         f_reg(31) <= "00000000000011101100011011000011";
         f_reg(32) <= "00000000010101011100100000000110";
         f_reg(33) <= "00000010100001011101000000100011";
         f_reg(34) <= "00111001110110111101011111110100";
         f_reg(35) <= "00000000000000000000000000000000";
         f_reg(36) <= "00000000010100101110000000101010";
         f_reg(37) <= "10101100000110100000001110110100";
         f_reg(38) <= "00000010101101101110100000100000";
         f_reg(39) <= "00000010001010001111000000100110";
         f_reg(40) <= "00000010000110010101000000100101";
         f_reg(41) <= "00000011100110000001100000100001";
         f_reg(42) <= "00000000011010100010000000100000";
         f_reg(43) <= "00000000000101000011001110000000";
         f_reg(44) <= "00000010110110000000100000100100";
         f_reg(45) <= "00000001111111010101100000100110";
         f_reg(46) <= "00000000000000000000000000000000";
         f_reg(47) <= "00111100000011011000001101011100";
         f_reg(48) <= "00000010111110011001100000100100";
         f_reg(49) <= "00000001010110000011100000100010";
         f_reg(50) <= "00000001100001100100100000000111";
         f_reg(51) <= "00000001001001000010100000100011";
         f_reg(52) <= "10101100000110110000001110111000";
         f_reg(53) <= "00000000111100110111000000100101";
         f_reg(54) <= "10101100000011100000001110111100";
         f_reg(55) <= "00000000000001010001000001000000";
         f_reg(56) <= "00110011110100101010011101011010";
         f_reg(57) <= "00000001011000101101000000000111";
         f_reg(58) <= "00000000000000011010110111000000";
         f_reg(59) <= "00000011101110001000100000101011";
         f_reg(60) <= "00000010101110100100000000000110";
         f_reg(61) <= "00100101101100000110000001101101";
         f_reg(62) <= "00000000000000000000000000000000";
         f_reg(63) <= "00000000000000000000000000000000";
         f_reg(64) <= "00000000000000000000000000000000";
         f_reg(65) <= "00000000000000000000000000000000";
         f_reg(66) <= "10101100000100000000001111000000";
         f_reg(67) <= "10101100000100010000001111000100";
         f_reg(68) <= "10101100000111010000001111001000";
         f_reg(69) <= "10101100000010000000001111001100";
         f_reg(70) <= "10101100000100100000001111010000";
         f_reg(71) <= "00100011111111111111111111111111";
         f_reg(72) <= "00011111111000001111111110111011";
         f_reg(73) <= "00010000000000000000000110100111";
         f_reg(74) <= "00111100000111100000001111100111";
         f_reg(75) <= "00111100000111110000001111100111";
         f_reg(76) <= "00000000000111101111010000000010";
         f_reg(77) <= "00000000000111111111110000000010";
         f_reg(78) <= "00111100000000010011010011001001";
         f_reg(79) <= "00111100000011110011010011001001";
         f_reg(80) <= "00111100000000101001011011000110";
         f_reg(81) <= "00111100000100001001011011000110";
         f_reg(82) <= "00000000000000010001100000000110";
         f_reg(83) <= "00000000000011111000100000000110";
         f_reg(84) <= "00101000001001000101110010010011";
         f_reg(85) <= "00101001111100100101110010010011";
         f_reg(86) <= "00010100100100100000000100001101";
         f_reg(87) <= "10101100000001000000001110101000";
         f_reg(88) <= "00000000000000000010100000100100";
         f_reg(89) <= "00000000000000001001100000100100";
         f_reg(90) <= "00000000001000000011000000000110";
         f_reg(91) <= "00000001111000001010000000000110";
         f_reg(92) <= "00000000110000010011100000100101";
         f_reg(93) <= "00000010100011111010100000100101";
         f_reg(94) <= "00000000000000000000000000000000";
         f_reg(95) <= "00000000000000000000000000000000";
         f_reg(96) <= "00000000110000000100000000100010";
         f_reg(97) <= "00000010100000001011000000100010";
         f_reg(98) <= "00000000000010000100110101000000";
         f_reg(99) <= "00000000000101101011110101000000";
         f_reg(100) <= "00100100101010101101000010011100";
         f_reg(101) <= "00100110011110001101000010011100";
         f_reg(102) <= "00000001010001010101100000100011";
         f_reg(103) <= "00000011000100111100100000100011";
         f_reg(104) <= "00101001011011000011010101010101";
         f_reg(105) <= "00101011001110100011010101010101";
         f_reg(106) <= "00000000011001000110100000100110";
         f_reg(107) <= "00000010001100101101100000100110";
         f_reg(108) <= "00000001100001100111000000101010";
         f_reg(109) <= "00000011010101001110000000101010";
         f_reg(110) <= "00101001110010101011100100100011";
         f_reg(111) <= "00101011100110001011100100100011";
         f_reg(112) <= "00000000001010110001100000000111";
         f_reg(113) <= "00000001111110011000100000000111";
         f_reg(114) <= "00010101000101100000000011110001";
         f_reg(115) <= "10101100000010000000001110101100";
         f_reg(116) <= "00000001101001110010000000000100";
         f_reg(117) <= "00000011011101011001000000000100";
         f_reg(118) <= "00000000000000000000000000000000";
         f_reg(119) <= "00000000000000000000000000000000";
         f_reg(120) <= "00000000010000010011000000100101";
         f_reg(121) <= "00000010000011111010000000100101";
         f_reg(122) <= "00000001011011000000100000100010";
         f_reg(123) <= "00000011001110100111100000100010";
         f_reg(124) <= "00010100010100000000000011100111";
         f_reg(125) <= "10101100000000100000001110110000";
         f_reg(126) <= "00000001100011010101100000100101";
         f_reg(127) <= "00000011010110111100100000100101";
         f_reg(128) <= "00000000000000010110111101000010";
         f_reg(129) <= "00000000000011111101111101000010";
         f_reg(130) <= "00000000110001110000100000100100";
         f_reg(131) <= "00000010100101010111100000100100";
         f_reg(132) <= "00110001001001110111010101110011";
         f_reg(133) <= "00110010111101010111010101110011";
         f_reg(134) <= "00000000000011100100111011000011";
         f_reg(135) <= "00000000000111001011111011000011";
         f_reg(136) <= "00010101001101110000000011011011";
         f_reg(137) <= "10101100000010010000001111010100";
         f_reg(138) <= "00000000010011010100100000000110";
         f_reg(139) <= "00000010000110111011100000000110";
         f_reg(140) <= "00010101100110100000000011010111";
         f_reg(141) <= "10101100000011000000001111011000";
         f_reg(142) <= "00000001011001010110000000100011";
         f_reg(143) <= "00000011001100111101000000100011";
         f_reg(144) <= "00111001110001011101011111110100";
         f_reg(145) <= "00111011100100111101011111110100";
         f_reg(146) <= "00000000000000000000000000000000";
         f_reg(147) <= "00000000000000000000000000000000";
         f_reg(148) <= "00000000010001100111000000101010";
         f_reg(149) <= "00000010000101001110000000101010";
         f_reg(150) <= "00010101100110100000000011001101";
         f_reg(151) <= "10101100000011000000001110110100";
         f_reg(152) <= "00000001101000010001000000100000";
         f_reg(153) <= "00000011011011111000000000100000";
         f_reg(154) <= "00000000100010000011000000100110";
         f_reg(155) <= "00000010010101101010000000100110";
         f_reg(156) <= "00000000011010010110000000100101";
         f_reg(157) <= "00000010001101111101000000100101";
         f_reg(158) <= "10001100000011010000001111010100";
         f_reg(159) <= "10001100000110110000001111010100";
         f_reg(160) <= "00010101101110111111111111111110";
         f_reg(161) <= "00000001110011010010000000100001";
         f_reg(162) <= "00000011100110111001000000100001";
         f_reg(163) <= "00000000100011000100000000100000";
         f_reg(164) <= "00000010010110101011000000100000";
         f_reg(165) <= "00000000000010110001101110000000";
         f_reg(166) <= "00000000000110011000101110000000";
         f_reg(167) <= "00000000001011010111000000100100";
         f_reg(168) <= "00000001111110111110000000100100";
         f_reg(169) <= "00000001010000100010000000100110";
         f_reg(170) <= "00000011000100001001000000100110";
         f_reg(171) <= "00000000000000000000000000000000";
         f_reg(172) <= "00000000000000000000000000000000";
         f_reg(173) <= "00111100000010111000001101011100";
         f_reg(174) <= "00111100000110011000001101011100";
         f_reg(175) <= "00000000111010010000100000100100";
         f_reg(176) <= "00000010101101110111100000100100";
         f_reg(177) <= "00000001100011010101000000100010";
         f_reg(178) <= "00000011010110111100000000100010";
         f_reg(179) <= "10001100000001110000001111011000";
         f_reg(180) <= "10001100000101010000001111011000";
         f_reg(181) <= "00010100111101011111111111111110";
         f_reg(182) <= "00000000111000110100100000000111";
         f_reg(183) <= "00000010101100011011100000000111";
         f_reg(184) <= "00000001001010000110000000100011";
         f_reg(185) <= "00000010111101101101000000100011";
         f_reg(186) <= "00010100101100110000000010101001";
         f_reg(187) <= "10101100000001010000001110111000";
         f_reg(188) <= "00000001010000010001100000100101";
         f_reg(189) <= "00000011000011111000100000100101";
         f_reg(190) <= "00010100011100010000000010100101";
         f_reg(191) <= "10101100000000110000001110111100";
         f_reg(192) <= "00000000000011000011100001000000";
         f_reg(193) <= "00000000000110101010100001000000";
         f_reg(194) <= "00110000110010011010011101011010";
         f_reg(195) <= "00110010100101111010011101011010";
         f_reg(196) <= "00000000100001110100000000000111";
         f_reg(197) <= "00000010010101011011000000000111";
         f_reg(198) <= "00000000000011100010110111000000";
         f_reg(199) <= "00000000000111001001110111000000";
         f_reg(200) <= "00000000010011010101000000101011";
         f_reg(201) <= "00000010000110111100000000101011";
         f_reg(202) <= "00000000101010000000100000000110";
         f_reg(203) <= "00000010011101100111100000000110";
         f_reg(204) <= "00100101011000110110000001101101";
         f_reg(205) <= "00100111001100010110000001101101";
         f_reg(206) <= "00000000000000000000000000000000";
         f_reg(207) <= "00000000000000000000000000000000";
         f_reg(208) <= "00000000000000000000000000000000";
         f_reg(209) <= "00000000000000000000000000000000";
         f_reg(210) <= "00000000000000000000000000000000";
         f_reg(211) <= "00000000000000000000000000000000";
         f_reg(212) <= "00000000000000000000000000000000";
         f_reg(213) <= "00000000000000000000000000000000";
         f_reg(214) <= "00010100011100010000000010001101";
         f_reg(215) <= "10101100000000110000001111000000";
         f_reg(216) <= "00010101010110000000000010001011";
         f_reg(217) <= "10101100000010100000001111000100";
         f_reg(218) <= "00010100010100000000000010001001";
         f_reg(219) <= "10101100000000100000001111001000";
         f_reg(220) <= "00010100001011110000000010000111";
         f_reg(221) <= "10101100000000010000001111001100";
         f_reg(222) <= "00010101001101110000000010000101";
         f_reg(223) <= "10101100000010010000001111010000";
         f_reg(224) <= "00100011110111011111111100000110";
         f_reg(225) <= "00010011101000000000000000010111";
         f_reg(226) <= "00100011110111011111111000001100";
         f_reg(227) <= "00010011101000000000000000010101";
         f_reg(228) <= "00100011110111011111110100010010";
         f_reg(229) <= "00010011101000000000000000010011";
         f_reg(230) <= "00100011110111101111111111111111";
         f_reg(231) <= "00100011111111111111111111111111";
         f_reg(232) <= "00010111110111110000000001111011";
         f_reg(233) <= "00011111111000001111111101100101";
         f_reg(234) <= "00010000000000000000000100000110";
         f_reg(235) <= "00000000000000000000000000000000";
         f_reg(236) <= "00000000000000000000000000000000";
         f_reg(237) <= "00000000000000000000000000000000";
         f_reg(238) <= "00000000000000000000000000000000";
         f_reg(239) <= "00000000000000000000000000000000";
         f_reg(240) <= "00000000000000000000000000000000";
         f_reg(241) <= "00000000000000000000000000000000";
         f_reg(242) <= "00000000000000000000000000000000";
         f_reg(243) <= "00000000000000000000000000000000";
         f_reg(244) <= "00000000000000000000000000000000";
         f_reg(245) <= "00000000000000000000000000000000";
         f_reg(246) <= "00000000000000000000000000000000";
         f_reg(247) <= "00000000000000000000000000000000";
         f_reg(248) <= "10001100000111010000011100110000";
         f_reg(249) <= "00011111101000000000000000000011";
         f_reg(250) <= "00100000000111010000000000111100";
         f_reg(251) <= "00010000000000000000000000000010";
         f_reg(252) <= "00100000000111010000000000000000";
         f_reg(253) <= "00010100001011110000000001100110";
         f_reg(254) <= "10101111101000010000011010111000";
         f_reg(255) <= "10001100000111010000011100110000";
         f_reg(256) <= "00011111101000000000000000000011";
         f_reg(257) <= "00100000000111010000000000111100";
         f_reg(258) <= "00010000000000000000000000000010";
         f_reg(259) <= "00100000000111010000000000000000";
         f_reg(260) <= "00010100010100000000000001011111";
         f_reg(261) <= "10101111101000100000011010111100";
         f_reg(262) <= "10001100000111010000011100110000";
         f_reg(263) <= "00011111101000000000000000000011";
         f_reg(264) <= "00100000000111010000000000111100";
         f_reg(265) <= "00010000000000000000000000000010";
         f_reg(266) <= "00100000000111010000000000000000";
         f_reg(267) <= "00010100011100010000000001011000";
         f_reg(268) <= "10101111101000110000011011000000";
         f_reg(269) <= "10001100000111010000011100110000";
         f_reg(270) <= "00011111101000000000000000000011";
         f_reg(271) <= "00100000000111010000000000111100";
         f_reg(272) <= "00010000000000000000000000000010";
         f_reg(273) <= "00100000000111010000000000000000";
         f_reg(274) <= "00010100100100100000000001010001";
         f_reg(275) <= "10101111101001000000011011000100";
         f_reg(276) <= "10001100000111010000011100110000";
         f_reg(277) <= "00011111101000000000000000000011";
         f_reg(278) <= "00100000000111010000000000111100";
         f_reg(279) <= "00010000000000000000000000000010";
         f_reg(280) <= "00100000000111010000000000000000";
         f_reg(281) <= "00010100101100110000000001001010";
         f_reg(282) <= "10101111101001010000011011001000";
         f_reg(283) <= "10001100000111010000011100110000";
         f_reg(284) <= "00011111101000000000000000000011";
         f_reg(285) <= "00100000000111010000000000111100";
         f_reg(286) <= "00010000000000000000000000000010";
         f_reg(287) <= "00100000000111010000000000000000";
         f_reg(288) <= "00010100110101000000000001000011";
         f_reg(289) <= "10101111101001100000011011001100";
         f_reg(290) <= "10001100000111010000011100110000";
         f_reg(291) <= "00011111101000000000000000000011";
         f_reg(292) <= "00100000000111010000000000111100";
         f_reg(293) <= "00010000000000000000000000000010";
         f_reg(294) <= "00100000000111010000000000000000";
         f_reg(295) <= "00010100111101010000000000111100";
         f_reg(296) <= "10101111101001110000011011010000";
         f_reg(297) <= "10001100000111010000011100110000";
         f_reg(298) <= "00011111101000000000000000000011";
         f_reg(299) <= "00100000000111010000000000111100";
         f_reg(300) <= "00010000000000000000000000000010";
         f_reg(301) <= "00100000000111010000000000000000";
         f_reg(302) <= "00010101000101100000000000110101";
         f_reg(303) <= "10101111101010000000011011010100";
         f_reg(304) <= "10001100000111010000011100110000";
         f_reg(305) <= "00011111101000000000000000000011";
         f_reg(306) <= "00100000000111010000000000111100";
         f_reg(307) <= "00010000000000000000000000000010";
         f_reg(308) <= "00100000000111010000000000000000";
         f_reg(309) <= "00010101001101110000000000101110";
         f_reg(310) <= "10101111101010010000011011011000";
         f_reg(311) <= "10001100000111010000011100110000";
         f_reg(312) <= "00011111101000000000000000000011";
         f_reg(313) <= "00100000000111010000000000111100";
         f_reg(314) <= "00010000000000000000000000000010";
         f_reg(315) <= "00100000000111010000000000000000";
         f_reg(316) <= "00010101010110000000000000100111";
         f_reg(317) <= "10101111101010100000011011011100";
         f_reg(318) <= "10001100000111010000011100110000";
         f_reg(319) <= "00011111101000000000000000000011";
         f_reg(320) <= "00100000000111010000000000111100";
         f_reg(321) <= "00010000000000000000000000000010";
         f_reg(322) <= "00100000000111010000000000000000";
         f_reg(323) <= "00010101011110010000000000100000";
         f_reg(324) <= "10101111101010110000011011100000";
         f_reg(325) <= "10001100000111010000011100110000";
         f_reg(326) <= "00011111101000000000000000000011";
         f_reg(327) <= "00100000000111010000000000111100";
         f_reg(328) <= "00010000000000000000000000000010";
         f_reg(329) <= "00100000000111010000000000000000";
         f_reg(330) <= "00010101100110100000000000011001";
         f_reg(331) <= "10101111101011000000011011100100";
         f_reg(332) <= "10001100000111010000011100110000";
         f_reg(333) <= "00011111101000000000000000000011";
         f_reg(334) <= "00100000000111010000000000111100";
         f_reg(335) <= "00010000000000000000000000000010";
         f_reg(336) <= "00100000000111010000000000000000";
         f_reg(337) <= "00010101101110110000000000010010";
         f_reg(338) <= "10101111101011010000011011101000";
         f_reg(339) <= "10001100000111010000011100110000";
         f_reg(340) <= "00011111101000000000000000000011";
         f_reg(341) <= "00100000000111010000000000111100";
         f_reg(342) <= "00010000000000000000000000000010";
         f_reg(343) <= "00100000000111010000000000000000";
         f_reg(344) <= "00010101110111000000000000001011";
         f_reg(345) <= "10101111101011100000011011101100";
         f_reg(346) <= "10001100000111010000011100110000";
         f_reg(347) <= "00011111101000000000000000000011";
         f_reg(348) <= "00100000000111010000000000111100";
         f_reg(349) <= "00010000000000000000000000000010";
         f_reg(350) <= "00100000000111010000000000000000";
         f_reg(351) <= "00010111110111110000000000000100";
         f_reg(352) <= "10101111101111100000011011110000";
         f_reg(353) <= "10101100000111010000011100110000";
         f_reg(354) <= "00010000000000001111111110000100";
         f_reg(355) <= "10001100000111010000011100110000";
         f_reg(356) <= "10001111101000010000011010111000";
         f_reg(357) <= "10001100000111010000011100110000";
         f_reg(358) <= "10001111101011110000011010111000";
         f_reg(359) <= "00010100001011111111111111111100";
         f_reg(360) <= "10001100000111010000011100110000";
         f_reg(361) <= "10001111101000100000011010111100";
         f_reg(362) <= "10001100000111010000011100110000";
         f_reg(363) <= "10001111101100000000011010111100";
         f_reg(364) <= "00010100010100001111111111111100";
         f_reg(365) <= "10001100000111010000011100110000";
         f_reg(366) <= "10001111101000110000011011000000";
         f_reg(367) <= "10001100000111010000011100110000";
         f_reg(368) <= "10001111101100010000011011000000";
         f_reg(369) <= "00010100011100011111111111111100";
         f_reg(370) <= "10001100000111010000011100110000";
         f_reg(371) <= "10001111101001000000011011000100";
         f_reg(372) <= "10001100000111010000011100110000";
         f_reg(373) <= "10001111101100100000011011000100";
         f_reg(374) <= "00010100100100101111111111111100";
         f_reg(375) <= "10001100000111010000011100110000";
         f_reg(376) <= "10001111101001010000011011001000";
         f_reg(377) <= "10001100000111010000011100110000";
         f_reg(378) <= "10001111101100110000011011001000";
         f_reg(379) <= "00010100101100111111111111111100";
         f_reg(380) <= "10001100000111010000011100110000";
         f_reg(381) <= "10001111101001100000011011001100";
         f_reg(382) <= "10001100000111010000011100110000";
         f_reg(383) <= "10001111101101000000011011001100";
         f_reg(384) <= "00010100110101001111111111111100";
         f_reg(385) <= "10001100000111010000011100110000";
         f_reg(386) <= "10001111101001110000011011010000";
         f_reg(387) <= "10001100000111010000011100110000";
         f_reg(388) <= "10001111101101010000011011010000";
         f_reg(389) <= "00010100111101011111111111111100";
         f_reg(390) <= "10001100000111010000011100110000";
         f_reg(391) <= "10001111101010000000011011010100";
         f_reg(392) <= "10001100000111010000011100110000";
         f_reg(393) <= "10001111101101100000011011010100";
         f_reg(394) <= "00010101000101101111111111111100";
         f_reg(395) <= "10001100000111010000011100110000";
         f_reg(396) <= "10001111101010010000011011011000";
         f_reg(397) <= "10001100000111010000011100110000";
         f_reg(398) <= "10001111101101110000011011011000";
         f_reg(399) <= "00010101001101111111111111111100";
         f_reg(400) <= "10001100000111010000011100110000";
         f_reg(401) <= "10001111101010100000011011011100";
         f_reg(402) <= "10001100000111010000011100110000";
         f_reg(403) <= "10001111101110000000011011011100";
         f_reg(404) <= "00010101010110001111111111111100";
         f_reg(405) <= "10001100000111010000011100110000";
         f_reg(406) <= "10001111101010110000011011100000";
         f_reg(407) <= "10001100000111010000011100110000";
         f_reg(408) <= "10001111101110010000011011100000";
         f_reg(409) <= "00010101011110011111111111111100";
         f_reg(410) <= "10001100000111010000011100110000";
         f_reg(411) <= "10001111101011000000011011100100";
         f_reg(412) <= "10001100000111010000011100110000";
         f_reg(413) <= "10001111101110100000011011100100";
         f_reg(414) <= "00010101100110101111111111111100";
         f_reg(415) <= "10001100000111010000011100110000";
         f_reg(416) <= "10001111101011010000011011101000";
         f_reg(417) <= "10001100000111010000011100110000";
         f_reg(418) <= "10001111101110110000011011101000";
         f_reg(419) <= "00010101101110111111111111111100";
         f_reg(420) <= "10001100000111010000011100110000";
         f_reg(421) <= "10001111101011100000011011101100";
         f_reg(422) <= "10001100000111010000011100110000";
         f_reg(423) <= "10001111101111000000011011101100";
         f_reg(424) <= "00010101110111001111111111111100";
         f_reg(425) <= "10001100000111010000011100110000";
         f_reg(426) <= "10001111101111100000011011110000";
         f_reg(427) <= "10001100000111010000011100110000";
         f_reg(428) <= "10001111101111110000011011110000";
         f_reg(429) <= "00010111110111111111111111111100";
         f_reg(430) <= "00010000000000001111111100111000";
         f_reg(431) <= "00000000000000000000000000000000";
         f_reg(432) <= "00000000000000000000000000000000";
         f_reg(433) <= "00000000000000000000000000000000";
         f_reg(434) <= "00000000000000000000000000000000";
         f_reg(435) <= "00000000000000000000000000000000";
         f_reg(436) <= "00000000000000000000000000000000";
         f_reg(437) <= "00000000000000000000000000000000";
         f_reg(438) <= "00000000000000000000000000000000";
         f_reg(439) <= "00000000000000000000000000000000";
         f_reg(440) <= "00000000000000000000000000000000";
         f_reg(441) <= "00000000000000000000000000000000";
         f_reg(442) <= "00000000000000000000000000000000";
         f_reg(443) <= "00000000000000000000000000000000";
         f_reg(444) <= "00000000000000000000000000000000";
         f_reg(445) <= "00000000000000000000000000000000";
         f_reg(446) <= "00000000000000000000000000000000";
         f_reg(447) <= "00000000000000000000000000000000";
         f_reg(448) <= "00000000000000000000000000000000";
         f_reg(449) <= "00000000000000000000000000000000";
         f_reg(450) <= "00000000000000000000000000000000";
         f_reg(451) <= "00000000000000000000000000000000";
         f_reg(452) <= "00000000000000000000000000000000";
         f_reg(453) <= "00000000000000000000000000000000";
         f_reg(454) <= "00000000000000000000000000000000";
         f_reg(455) <= "00000000000000000000000000000000";
         f_reg(456) <= "00000000000000000000000000000000";
         f_reg(457) <= "00000000000000000000000000000000";
         f_reg(458) <= "00000000000000000000000000000000";
         f_reg(459) <= "00000000000000000000000000000000";
         f_reg(460) <= "00000000000000000000000000000000";
         f_reg(461) <= "00000000000000000000001111100111";
         f_reg(462) <= "00000000000000000000000000000000";
         f_reg(463) <= "00000000000000000000000000000000";
         f_reg(464) <= "00000000000000000000000000000000";
         f_reg(465) <= "00000000000000000000000000000000";
         f_reg(466) <= "00000000000000000000000000000000";
         f_reg(467) <= "00000000000000000000000000000000";
         f_reg(468) <= "00000000000000000000000000000000";
         f_reg(469) <= "00000000000000000000000000000000";
         f_reg(470) <= "00000000000000000000000000000000";
         f_reg(471) <= "00000000000000000000000000000000";
         f_reg(472) <= "00000000000000000000000000000000";
         f_reg(473) <= "00000000000000000000000000000000";
         f_reg(474) <= "00000000000000000000000000000000";
         f_reg(475) <= "00000000000000000000000000000000";
         f_reg(476) <= "00000000000000000000000000000000";
         f_reg(477) <= "00000000000000000000000000000000";
         f_reg(478) <= "00000000000000000000000000000000";
         f_reg(479) <= "00000000000000000000000000000000";
         f_reg(480) <= "00000000000000000000000000000000";
         f_reg(481) <= "00000000000000000000000000000000";
         f_reg(482) <= "00000000000000000000000000000000";
         f_reg(483) <= "00000000000000000000000000000000";
         f_reg(484) <= "00000000000000000000000000000000";
         f_reg(485) <= "00000000000000000000000000000000";
         f_reg(486) <= "00000000000000000000000000000000";
         f_reg(487) <= "00000000000000000000000000000000";
         f_reg(488) <= "00000000000000000000000000000000";
         f_reg(489) <= "00000000000000000000000000000000";
         f_reg(490) <= "00000000000000000000000000000000";
         f_reg(491) <= "00000000000000000000000000000000";
         f_reg(492) <= "00000000000000000000000000000000";
         f_reg(493) <= "00000000000000000000000000000000";
         f_reg(494) <= "00000000000000000000000000000000";
         f_reg(495) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 13513
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- LUI R2 -26938
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SRLV R3 R1 R0
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SLTI R4 R1 23699
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SW R4 R0 936
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- AND R5 R0 R0
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- SRLV R6 R0 R1
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- OR R7 R6 R1
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- NOP
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- SUB R8 R6 R0
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- SLL R9 R8 21
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- ADDIU R10 R5 -12132
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- SUBU R11 R10 R5
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- SLTI R12 R11 13653
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- XOR R13 R3 R4
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- SLT R14 R12 R6
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SLTI R15 R14 -18141
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- SRAV R16 R11 R1
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SW R8 R0 940
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- SLLV R17 R7 R13
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- NOP
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- OR R18 R2 R1
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- SUB R19 R11 R12
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- SW R2 R0 944
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- OR R20 R12 R13
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- SRL R21 R19 29
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- AND R22 R18 R7
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- ANDI R23 R9 30067
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- SRA R24 R14 27
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- SRLV R25 R21 R2
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- SUBU R26 R20 R5
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- XORI R27 R14 -10252
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- NOP
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- SLT R28 R2 R18
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- SW R26 R0 948
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- ADD R29 R21 R22
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- XOR R30 R17 R8
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- OR R10 R16 R25
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- ADDU R3 R28 R24
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- ADD R4 R3 R10
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SLL R6 R20 14
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- AND R1 R22 R24
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- XOR R11 R15 R29
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- NOP
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- LUI R13 -31908
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- AND R19 R23 R25
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- SUB R7 R10 R24
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- SRAV R9 R6 R12
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SUBU R5 R9 R4
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- SW R27 R0 952
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- OR R14 R7 R19
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SW R14 R0 956
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SLL R2 R5 1
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- ANDI R18 R30 -22694
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SRAV R26 R2 R11
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- SLL R21 R1 23
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- SLTU R17 R29 R24
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SRLV R8 R26 R21
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- ADDIU R16 R13 24685
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- NOP
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- NOP
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- NOP
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- NOP
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- SW R16 R0 960
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- SW R17 R0 964
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- SW R29 R0 968
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- SW R8 R0 972
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SW R18 R0 976
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- BGTZ R31 -69
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- BEQ R0 R0 423
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- LUI R30 999
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- LUI R31 999
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- LUI R1 13513
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- LUI R15 13513
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- LUI R2 -26938
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- LUI R16 -26938
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- SRLV R3 R1 R0
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SRLV R17 R15 R0
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- SLTI R4 R1 23699
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- SLTI R18 R15 23699
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- BNE R4 R18 269
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SW R4 R0 936
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- AND R5 R0 R0
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- AND R19 R0 R0
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- SRLV R6 R0 R1
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- SRLV R20 R0 R15
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- OR R7 R6 R1
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- OR R21 R20 R15
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- NOP
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- NOP
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- SUB R8 R6 R0
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SUB R22 R20 R0
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SLL R9 R8 21
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- SLL R23 R22 21
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- ADDIU R10 R5 -12132
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- ADDIU R24 R19 -12132
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- SUBU R11 R10 R5
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SUBU R25 R24 R19
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- SLTI R12 R11 13653
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- SLTI R26 R25 13653
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- XOR R13 R3 R4
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- XOR R27 R17 R18
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- SLT R14 R12 R6
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- SLT R28 R26 R20
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- SLTI R10 R14 -18141
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- SLTI R24 R28 -18141
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- SRAV R3 R11 R1
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- SRAV R17 R25 R15
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- BNE R8 R22 241
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- SW R8 R0 940
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- SLLV R4 R7 R13
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- SLLV R18 R21 R27
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- NOP
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- NOP
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- OR R6 R2 R1
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- OR R20 R16 R15
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- SUB R1 R11 R12
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- SUB R15 R25 R26
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- BNE R2 R16 231
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- SW R2 R0 944
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- OR R11 R12 R13
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- OR R25 R26 R27
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SRL R13 R1 29
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- SRL R27 R15 29
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- AND R1 R6 R7
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- AND R15 R20 R21
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- ANDI R7 R9 30067
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- ANDI R21 R23 30067
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- SRA R9 R14 27
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- SRA R23 R28 27
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- BNE R9 R23 219
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- SW R9 R0 980
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SRLV R9 R13 R2
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- SRLV R23 R27 R16
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- BNE R12 R26 215
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- SW R12 R0 984
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- SUBU R12 R11 R5
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- SUBU R26 R25 R19
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- XORI R5 R14 -10252
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- XORI R19 R28 -10252
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- NOP
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- NOP
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- SLT R14 R2 R6
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- SLT R28 R16 R20
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- BNE R12 R26 205
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- SW R12 R0 948
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- ADD R2 R13 R1
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- ADD R16 R27 R15
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- XOR R6 R4 R8
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- XOR R20 R18 R22
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- OR R12 R3 R9
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- OR R26 R17 R23
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- LW R13 R0 980
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- LW R27 R0 980
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- BNE R13 R27 -2
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- ADDU R4 R14 R13
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- ADDU R18 R28 R27
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- ADD R8 R4 R12
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- ADD R22 R18 R26
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- SLL R3 R11 14
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- SLL R17 R25 14
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- AND R14 R1 R13
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- AND R28 R15 R27
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- XOR R4 R10 R2
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- XOR R18 R24 R16
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- NOP
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- NOP
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- LUI R11 -31908
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- LUI R25 -31908
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- AND R1 R7 R9
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- AND R15 R21 R23
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- SUB R10 R12 R13
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- SUB R24 R26 R27
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- LW R7 R0 984
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- LW R21 R0 984
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- BNE R7 R21 -2
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SRAV R9 R3 R7
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- SRAV R23 R17 R21
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- SUBU R12 R9 R8
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- SUBU R26 R23 R22
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- BNE R5 R19 169
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- SW R5 R0 952
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- OR R3 R10 R1
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- OR R17 R24 R15
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- BNE R3 R17 165
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- SW R3 R0 956
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- SLL R7 R12 1
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- SLL R21 R26 1
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- ANDI R9 R6 -22694
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- ANDI R23 R20 -22694
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- SRAV R8 R7 R4
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- SRAV R22 R21 R18
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- SLL R5 R14 23
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- SLL R19 R28 23
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- SLTU R10 R2 R13
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- SLTU R24 R16 R27
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- SRLV R1 R8 R5
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- SRLV R15 R22 R19
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- ADDIU R3 R11 24685
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- ADDIU R17 R25 24685
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- NOP
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- NOP
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- NOP
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- NOP
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- NOP
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- NOP
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- NOP
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- NOP
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- BNE R3 R17 141
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- SW R3 R0 960
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- BNE R10 R24 139
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- SW R10 R0 964
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- BNE R2 R16 137
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- SW R2 R0 968
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- BNE R1 R15 135
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- SW R1 R0 972
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- BNE R9 R23 133
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- SW R9 R0 976
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- BEQ R29 R0 23
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- BEQ R29 R0 21
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- BEQ R29 R0 19
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- BNE R30 R31 123
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- BGTZ R31 -155
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- BEQ R0 R0 262
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- NOP
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- NOP
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- NOP
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- NOP
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- NOP
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- NOP
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- NOP
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- NOP
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- NOP
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- NOP
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- NOP
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- NOP
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- NOP
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- SW R1 R29 1720
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- SW R2 R29 1724
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- SW R3 R29 1728
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- SW R4 R29 1732
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- SW R5 R29 1736
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- SW R6 R29 1740
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- SW R7 R29 1744
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- SW R8 R29 1748
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- SW R9 R29 1752
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- SW R10 R29 1756
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- SW R11 R29 1760
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- SW R12 R29 1764
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- SW R13 R29 1768
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- SW R14 R29 1772
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- SW R30 R29 1776
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- SW R29 R0 1840
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- BEQ R0 R0 -124
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- LW R1 R29 1720
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- LW R15 R29 1720
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- LW R2 R29 1724
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- LW R16 R29 1724
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- LW R3 R29 1728
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- LW R17 R29 1728
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- LW R4 R29 1732
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- LW R18 R29 1732
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- LW R5 R29 1736
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- LW R19 R29 1736
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- LW R6 R29 1740
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- LW R20 R29 1740
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- LW R7 R29 1744
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- LW R21 R29 1744
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- LW R8 R29 1748
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- LW R22 R29 1748
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- LW R9 R29 1752
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- LW R23 R29 1752
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- LW R10 R29 1756
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- LW R24 R29 1756
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- LW R11 R29 1760
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- LW R25 R29 1760
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- LW R12 R29 1764
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- LW R26 R29 1764
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- LW R13 R29 1768
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- LW R27 R29 1768
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- LW R14 R29 1772
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- LW R28 R29 1772
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R30 R29 1776
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- LW R29 R0 1840
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- LW R31 R29 1776
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- BEQ R0 R0 -200
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- NOP
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- NOP
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- NOP
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- NOP
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- NOP
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- NOP
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- NOP
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- NOP
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- NOP
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- NOP
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- NOP
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- NOP
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- NOP
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- NOP
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- NOP
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- NOP
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- NOP
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- NOP
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- NOP
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- NOP
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- NOP
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- NOP
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- NOP
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- NOP
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- NOP
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- NOP
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- NOP
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- NOP
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- NOP
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- NOP
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- NOP
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- NOP
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- NOP
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- NOP
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- NOP
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- NOP
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- NOP
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- NOP
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- NOP
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- NOP
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- NOP
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- NOP
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- NOP
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- NOP
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- NOP
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- NOP
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- NOP
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- NOP
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- NOP
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- NOP
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- NOP
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- NOP
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- NOP
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- NOP
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- NOP
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- NOP
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- NOP
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- NOP
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- NOP
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- NOP
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- NOP
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- NOP
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- NOP
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- NOP
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- NOP
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010011010011001001";
                        f_reg(4) <= "00111100000000101001011011000110";
                        f_reg(5) <= "00000000000000010001100000000110";
                        f_reg(6) <= "00101000001001000101110010010011";
                        f_reg(7) <= "10101100000001000000001110101000";
                        f_reg(8) <= "00000000000000000010100000100100";
                        f_reg(9) <= "00000000001000000011000000000110";
                        f_reg(10) <= "00000000110000010011100000100101";
                        f_reg(11) <= "00000000000000000000000000000000";
                        f_reg(12) <= "00000000110000000100000000100010";
                        f_reg(13) <= "00000000000010000100110101000000";
                        f_reg(14) <= "00100100101010101101000010011100";
                        f_reg(15) <= "00000001010001010101100000100011";
                        f_reg(16) <= "00101001011011000011010101010101";
                        f_reg(17) <= "00000000011001000110100000100110";
                        f_reg(18) <= "00000001100001100111000000101010";
                        f_reg(19) <= "00101001110011111011100100100011";
                        f_reg(20) <= "00000000001010111000000000000111";
                        f_reg(21) <= "10101100000010000000001110101100";
                        f_reg(22) <= "00000001101001111000100000000100";
                        f_reg(23) <= "00000000000000000000000000000000";
                        f_reg(24) <= "00000000010000011001000000100101";
                        f_reg(25) <= "00000001011011001001100000100010";
                        f_reg(26) <= "10101100000000100000001110110000";
                        f_reg(27) <= "00000001100011011010000000100101";
                        f_reg(28) <= "00000000000100111010111101000010";
                        f_reg(29) <= "00000010010001111011000000100100";
                        f_reg(30) <= "00110001001101110111010101110011";
                        f_reg(31) <= "00000000000011101100011011000011";
                        f_reg(32) <= "00000000010101011100100000000110";
                        f_reg(33) <= "00000010100001011101000000100011";
                        f_reg(34) <= "00111001110110111101011111110100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000000010100101110000000101010";
                        f_reg(37) <= "10101100000110100000001110110100";
                        f_reg(38) <= "00000010101101101110100000100000";
                        f_reg(39) <= "00000010001010001111000000100110";
                        f_reg(40) <= "00000010000110010101000000100101";
                        f_reg(41) <= "00000011100110000001100000100001";
                        f_reg(42) <= "00000000011010100010000000100000";
                        f_reg(43) <= "00000000000101000011001110000000";
                        f_reg(44) <= "00000010110110000000100000100100";
                        f_reg(45) <= "00000001111111010101100000100110";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00111100000011011000001101011100";
                        f_reg(48) <= "00000010111110011001100000100100";
                        f_reg(49) <= "00000001010110000011100000100010";
                        f_reg(50) <= "00000001100001100100100000000111";
                        f_reg(51) <= "00000001001001000010100000100011";
                        f_reg(52) <= "10101100000110110000001110111000";
                        f_reg(53) <= "00000000111100110111000000100101";
                        f_reg(54) <= "10101100000011100000001110111100";
                        f_reg(55) <= "00000000000001010001000001000000";
                        f_reg(56) <= "00110011110100101010011101011010";
                        f_reg(57) <= "00000001011000101101000000000111";
                        f_reg(58) <= "00000000000000011010110111000000";
                        f_reg(59) <= "00000011101110001000100000101011";
                        f_reg(60) <= "00000010101110100100000000000110";
                        f_reg(61) <= "00100101101100000110000001101101";
                        f_reg(62) <= "00000000000000000000000000000000";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000000000000000000000000000000";
                        f_reg(66) <= "10101100000100000000001111000000";
                        f_reg(67) <= "10101100000100010000001111000100";
                        f_reg(68) <= "10101100000111010000001111001000";
                        f_reg(69) <= "10101100000010000000001111001100";
                        f_reg(70) <= "10101100000100100000001111010000";
                        f_reg(71) <= "00100011111111111111111111111111";
                        f_reg(72) <= "00011111111000001111111110111011";
                        f_reg(73) <= "00010000000000000000000110100111";
                        f_reg(74) <= "00111100000111100000001111100111";
                        f_reg(75) <= "00111100000111110000001111100111";
                        f_reg(76) <= "00000000000111101111010000000010";
                        f_reg(77) <= "00000000000111111111110000000010";
                        f_reg(78) <= "00111100000000010011010011001001";
                        f_reg(79) <= "00111100000011110011010011001001";
                        f_reg(80) <= "00111100000000101001011011000110";
                        f_reg(81) <= "00111100000100001001011011000110";
                        f_reg(82) <= "00000000000000010001100000000110";
                        f_reg(83) <= "00000000000011111000100000000110";
                        f_reg(84) <= "00101000001001000101110010010011";
                        f_reg(85) <= "00101001111100100101110010010011";
                        f_reg(86) <= "00010100100100100000000100001101";
                        f_reg(87) <= "10101100000001000000001110101000";
                        f_reg(88) <= "00000000000000000010100000100100";
                        f_reg(89) <= "00000000000000001001100000100100";
                        f_reg(90) <= "00000000001000000011000000000110";
                        f_reg(91) <= "00000001111000001010000000000110";
                        f_reg(92) <= "00000000110000010011100000100101";
                        f_reg(93) <= "00000010100011111010100000100101";
                        f_reg(94) <= "00000000000000000000000000000000";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000110000000100000000100010";
                        f_reg(97) <= "00000010100000001011000000100010";
                        f_reg(98) <= "00000000000010000100110101000000";
                        f_reg(99) <= "00000000000101101011110101000000";
                        f_reg(100) <= "00100100101010101101000010011100";
                        f_reg(101) <= "00100110011110001101000010011100";
                        f_reg(102) <= "00000001010001010101100000100011";
                        f_reg(103) <= "00000011000100111100100000100011";
                        f_reg(104) <= "00101001011011000011010101010101";
                        f_reg(105) <= "00101011001110100011010101010101";
                        f_reg(106) <= "00000000011001000110100000100110";
                        f_reg(107) <= "00000010001100101101100000100110";
                        f_reg(108) <= "00000001100001100111000000101010";
                        f_reg(109) <= "00000011010101001110000000101010";
                        f_reg(110) <= "00101001110010101011100100100011";
                        f_reg(111) <= "00101011100110001011100100100011";
                        f_reg(112) <= "00000000001010110001100000000111";
                        f_reg(113) <= "00000001111110011000100000000111";
                        f_reg(114) <= "00010101000101100000000011110001";
                        f_reg(115) <= "10101100000010000000001110101100";
                        f_reg(116) <= "00000001101001110010000000000100";
                        f_reg(117) <= "00000011011101011001000000000100";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000010000010011000000100101";
                        f_reg(121) <= "00000010000011111010000000100101";
                        f_reg(122) <= "00000001011011000000100000100010";
                        f_reg(123) <= "00000011001110100111100000100010";
                        f_reg(124) <= "00010100010100000000000011100111";
                        f_reg(125) <= "10101100000000100000001110110000";
                        f_reg(126) <= "00000001100011010101100000100101";
                        f_reg(127) <= "00000011010110111100100000100101";
                        f_reg(128) <= "00000000000000010110111101000010";
                        f_reg(129) <= "00000000000011111101111101000010";
                        f_reg(130) <= "00000000110001110000100000100100";
                        f_reg(131) <= "00000010100101010111100000100100";
                        f_reg(132) <= "00110001001001110111010101110011";
                        f_reg(133) <= "00110010111101010111010101110011";
                        f_reg(134) <= "00000000000011100100111011000011";
                        f_reg(135) <= "00000000000111001011111011000011";
                        f_reg(136) <= "00010101001101110000000011011011";
                        f_reg(137) <= "10101100000010010000001111010100";
                        f_reg(138) <= "00000000010011010100100000000110";
                        f_reg(139) <= "00000010000110111011100000000110";
                        f_reg(140) <= "00010101100110100000000011010111";
                        f_reg(141) <= "10101100000011000000001111011000";
                        f_reg(142) <= "00000001011001010110000000100011";
                        f_reg(143) <= "00000011001100111101000000100011";
                        f_reg(144) <= "00111001110001011101011111110100";
                        f_reg(145) <= "00111011100100111101011111110100";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000010001100111000000101010";
                        f_reg(149) <= "00000010000101001110000000101010";
                        f_reg(150) <= "00010101100110100000000011001101";
                        f_reg(151) <= "10101100000011000000001110110100";
                        f_reg(152) <= "00000001101000010001000000100000";
                        f_reg(153) <= "00000011011011111000000000100000";
                        f_reg(154) <= "00000000100010000011000000100110";
                        f_reg(155) <= "00000010010101101010000000100110";
                        f_reg(156) <= "00000000011010010110000000100101";
                        f_reg(157) <= "00000010001101111101000000100101";
                        f_reg(158) <= "10001100000011010000001111010100";
                        f_reg(159) <= "10001100000110110000001111010100";
                        f_reg(160) <= "00010101101110111111111111111110";
                        f_reg(161) <= "00000001110011010010000000100001";
                        f_reg(162) <= "00000011100110111001000000100001";
                        f_reg(163) <= "00000000100011000100000000100000";
                        f_reg(164) <= "00000010010110101011000000100000";
                        f_reg(165) <= "00000000000010110001101110000000";
                        f_reg(166) <= "00000000000110011000101110000000";
                        f_reg(167) <= "00000000001011010111000000100100";
                        f_reg(168) <= "00000001111110111110000000100100";
                        f_reg(169) <= "00000001010000100010000000100110";
                        f_reg(170) <= "00000011000100001001000000100110";
                        f_reg(171) <= "00000000000000000000000000000000";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00111100000010111000001101011100";
                        f_reg(174) <= "00111100000110011000001101011100";
                        f_reg(175) <= "00000000111010010000100000100100";
                        f_reg(176) <= "00000010101101110111100000100100";
                        f_reg(177) <= "00000001100011010101000000100010";
                        f_reg(178) <= "00000011010110111100000000100010";
                        f_reg(179) <= "10001100000001110000001111011000";
                        f_reg(180) <= "10001100000101010000001111011000";
                        f_reg(181) <= "00010100111101011111111111111110";
                        f_reg(182) <= "00000000111000110100100000000111";
                        f_reg(183) <= "00000010101100011011100000000111";
                        f_reg(184) <= "00000001001010000110000000100011";
                        f_reg(185) <= "00000010111101101101000000100011";
                        f_reg(186) <= "00010100101100110000000010101001";
                        f_reg(187) <= "10101100000001010000001110111000";
                        f_reg(188) <= "00000001010000010001100000100101";
                        f_reg(189) <= "00000011000011111000100000100101";
                        f_reg(190) <= "00010100011100010000000010100101";
                        f_reg(191) <= "10101100000000110000001110111100";
                        f_reg(192) <= "00000000000011000011100001000000";
                        f_reg(193) <= "00000000000110101010100001000000";
                        f_reg(194) <= "00110000110010011010011101011010";
                        f_reg(195) <= "00110010100101111010011101011010";
                        f_reg(196) <= "00000000100001110100000000000111";
                        f_reg(197) <= "00000010010101011011000000000111";
                        f_reg(198) <= "00000000000011100010110111000000";
                        f_reg(199) <= "00000000000111001001110111000000";
                        f_reg(200) <= "00000000010011010101000000101011";
                        f_reg(201) <= "00000010000110111100000000101011";
                        f_reg(202) <= "00000000101010000000100000000110";
                        f_reg(203) <= "00000010011101100111100000000110";
                        f_reg(204) <= "00100101011000110110000001101101";
                        f_reg(205) <= "00100111001100010110000001101101";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00010100011100010000000010001101";
                        f_reg(215) <= "10101100000000110000001111000000";
                        f_reg(216) <= "00010101010110000000000010001011";
                        f_reg(217) <= "10101100000010100000001111000100";
                        f_reg(218) <= "00010100010100000000000010001001";
                        f_reg(219) <= "10101100000000100000001111001000";
                        f_reg(220) <= "00010100001011110000000010000111";
                        f_reg(221) <= "10101100000000010000001111001100";
                        f_reg(222) <= "00010101001101110000000010000101";
                        f_reg(223) <= "10101100000010010000001111010000";
                        f_reg(224) <= "00100011110111011111111100000110";
                        f_reg(225) <= "00010011101000000000000000010111";
                        f_reg(226) <= "00100011110111011111111000001100";
                        f_reg(227) <= "00010011101000000000000000010101";
                        f_reg(228) <= "00100011110111011111110100010010";
                        f_reg(229) <= "00010011101000000000000000010011";
                        f_reg(230) <= "00100011110111101111111111111111";
                        f_reg(231) <= "00100011111111111111111111111111";
                        f_reg(232) <= "00010111110111110000000001111011";
                        f_reg(233) <= "00011111111000001111111101100101";
                        f_reg(234) <= "00010000000000000000000100000110";
                        f_reg(235) <= "00000000000000000000000000000000";
                        f_reg(236) <= "00000000000000000000000000000000";
                        f_reg(237) <= "00000000000000000000000000000000";
                        f_reg(238) <= "00000000000000000000000000000000";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000000000000000000000000000000";
                        f_reg(242) <= "00000000000000000000000000000000";
                        f_reg(243) <= "00000000000000000000000000000000";
                        f_reg(244) <= "00000000000000000000000000000000";
                        f_reg(245) <= "00000000000000000000000000000000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "10001100000111010000011100110000";
                        f_reg(249) <= "00011111101000000000000000000011";
                        f_reg(250) <= "00100000000111010000000000111100";
                        f_reg(251) <= "00010000000000000000000000000010";
                        f_reg(252) <= "00100000000111010000000000000000";
                        f_reg(253) <= "00010100001011110000000001100110";
                        f_reg(254) <= "10101111101000010000011010111000";
                        f_reg(255) <= "10001100000111010000011100110000";
                        f_reg(256) <= "00011111101000000000000000000011";
                        f_reg(257) <= "00100000000111010000000000111100";
                        f_reg(258) <= "00010000000000000000000000000010";
                        f_reg(259) <= "00100000000111010000000000000000";
                        f_reg(260) <= "00010100010100000000000001011111";
                        f_reg(261) <= "10101111101000100000011010111100";
                        f_reg(262) <= "10001100000111010000011100110000";
                        f_reg(263) <= "00011111101000000000000000000011";
                        f_reg(264) <= "00100000000111010000000000111100";
                        f_reg(265) <= "00010000000000000000000000000010";
                        f_reg(266) <= "00100000000111010000000000000000";
                        f_reg(267) <= "00010100011100010000000001011000";
                        f_reg(268) <= "10101111101000110000011011000000";
                        f_reg(269) <= "10001100000111010000011100110000";
                        f_reg(270) <= "00011111101000000000000000000011";
                        f_reg(271) <= "00100000000111010000000000111100";
                        f_reg(272) <= "00010000000000000000000000000010";
                        f_reg(273) <= "00100000000111010000000000000000";
                        f_reg(274) <= "00010100100100100000000001010001";
                        f_reg(275) <= "10101111101001000000011011000100";
                        f_reg(276) <= "10001100000111010000011100110000";
                        f_reg(277) <= "00011111101000000000000000000011";
                        f_reg(278) <= "00100000000111010000000000111100";
                        f_reg(279) <= "00010000000000000000000000000010";
                        f_reg(280) <= "00100000000111010000000000000000";
                        f_reg(281) <= "00010100101100110000000001001010";
                        f_reg(282) <= "10101111101001010000011011001000";
                        f_reg(283) <= "10001100000111010000011100110000";
                        f_reg(284) <= "00011111101000000000000000000011";
                        f_reg(285) <= "00100000000111010000000000111100";
                        f_reg(286) <= "00010000000000000000000000000010";
                        f_reg(287) <= "00100000000111010000000000000000";
                        f_reg(288) <= "00010100110101000000000001000011";
                        f_reg(289) <= "10101111101001100000011011001100";
                        f_reg(290) <= "10001100000111010000011100110000";
                        f_reg(291) <= "00011111101000000000000000000011";
                        f_reg(292) <= "00100000000111010000000000111100";
                        f_reg(293) <= "00010000000000000000000000000010";
                        f_reg(294) <= "00100000000111010000000000000000";
                        f_reg(295) <= "00010100111101010000000000111100";
                        f_reg(296) <= "10101111101001110000011011010000";
                        f_reg(297) <= "10001100000111010000011100110000";
                        f_reg(298) <= "00011111101000000000000000000011";
                        f_reg(299) <= "00100000000111010000000000111100";
                        f_reg(300) <= "00010000000000000000000000000010";
                        f_reg(301) <= "00100000000111010000000000000000";
                        f_reg(302) <= "00010101000101100000000000110101";
                        f_reg(303) <= "10101111101010000000011011010100";
                        f_reg(304) <= "10001100000111010000011100110000";
                        f_reg(305) <= "00011111101000000000000000000011";
                        f_reg(306) <= "00100000000111010000000000111100";
                        f_reg(307) <= "00010000000000000000000000000010";
                        f_reg(308) <= "00100000000111010000000000000000";
                        f_reg(309) <= "00010101001101110000000000101110";
                        f_reg(310) <= "10101111101010010000011011011000";
                        f_reg(311) <= "10001100000111010000011100110000";
                        f_reg(312) <= "00011111101000000000000000000011";
                        f_reg(313) <= "00100000000111010000000000111100";
                        f_reg(314) <= "00010000000000000000000000000010";
                        f_reg(315) <= "00100000000111010000000000000000";
                        f_reg(316) <= "00010101010110000000000000100111";
                        f_reg(317) <= "10101111101010100000011011011100";
                        f_reg(318) <= "10001100000111010000011100110000";
                        f_reg(319) <= "00011111101000000000000000000011";
                        f_reg(320) <= "00100000000111010000000000111100";
                        f_reg(321) <= "00010000000000000000000000000010";
                        f_reg(322) <= "00100000000111010000000000000000";
                        f_reg(323) <= "00010101011110010000000000100000";
                        f_reg(324) <= "10101111101010110000011011100000";
                        f_reg(325) <= "10001100000111010000011100110000";
                        f_reg(326) <= "00011111101000000000000000000011";
                        f_reg(327) <= "00100000000111010000000000111100";
                        f_reg(328) <= "00010000000000000000000000000010";
                        f_reg(329) <= "00100000000111010000000000000000";
                        f_reg(330) <= "00010101100110100000000000011001";
                        f_reg(331) <= "10101111101011000000011011100100";
                        f_reg(332) <= "10001100000111010000011100110000";
                        f_reg(333) <= "00011111101000000000000000000011";
                        f_reg(334) <= "00100000000111010000000000111100";
                        f_reg(335) <= "00010000000000000000000000000010";
                        f_reg(336) <= "00100000000111010000000000000000";
                        f_reg(337) <= "00010101101110110000000000010010";
                        f_reg(338) <= "10101111101011010000011011101000";
                        f_reg(339) <= "10001100000111010000011100110000";
                        f_reg(340) <= "00011111101000000000000000000011";
                        f_reg(341) <= "00100000000111010000000000111100";
                        f_reg(342) <= "00010000000000000000000000000010";
                        f_reg(343) <= "00100000000111010000000000000000";
                        f_reg(344) <= "00010101110111000000000000001011";
                        f_reg(345) <= "10101111101011100000011011101100";
                        f_reg(346) <= "10001100000111010000011100110000";
                        f_reg(347) <= "00011111101000000000000000000011";
                        f_reg(348) <= "00100000000111010000000000111100";
                        f_reg(349) <= "00010000000000000000000000000010";
                        f_reg(350) <= "00100000000111010000000000000000";
                        f_reg(351) <= "00010111110111110000000000000100";
                        f_reg(352) <= "10101111101111100000011011110000";
                        f_reg(353) <= "10101100000111010000011100110000";
                        f_reg(354) <= "00010000000000001111111110000100";
                        f_reg(355) <= "10001100000111010000011100110000";
                        f_reg(356) <= "10001111101000010000011010111000";
                        f_reg(357) <= "10001100000111010000011100110000";
                        f_reg(358) <= "10001111101011110000011010111000";
                        f_reg(359) <= "00010100001011111111111111111100";
                        f_reg(360) <= "10001100000111010000011100110000";
                        f_reg(361) <= "10001111101000100000011010111100";
                        f_reg(362) <= "10001100000111010000011100110000";
                        f_reg(363) <= "10001111101100000000011010111100";
                        f_reg(364) <= "00010100010100001111111111111100";
                        f_reg(365) <= "10001100000111010000011100110000";
                        f_reg(366) <= "10001111101000110000011011000000";
                        f_reg(367) <= "10001100000111010000011100110000";
                        f_reg(368) <= "10001111101100010000011011000000";
                        f_reg(369) <= "00010100011100011111111111111100";
                        f_reg(370) <= "10001100000111010000011100110000";
                        f_reg(371) <= "10001111101001000000011011000100";
                        f_reg(372) <= "10001100000111010000011100110000";
                        f_reg(373) <= "10001111101100100000011011000100";
                        f_reg(374) <= "00010100100100101111111111111100";
                        f_reg(375) <= "10001100000111010000011100110000";
                        f_reg(376) <= "10001111101001010000011011001000";
                        f_reg(377) <= "10001100000111010000011100110000";
                        f_reg(378) <= "10001111101100110000011011001000";
                        f_reg(379) <= "00010100101100111111111111111100";
                        f_reg(380) <= "10001100000111010000011100110000";
                        f_reg(381) <= "10001111101001100000011011001100";
                        f_reg(382) <= "10001100000111010000011100110000";
                        f_reg(383) <= "10001111101101000000011011001100";
                        f_reg(384) <= "00010100110101001111111111111100";
                        f_reg(385) <= "10001100000111010000011100110000";
                        f_reg(386) <= "10001111101001110000011011010000";
                        f_reg(387) <= "10001100000111010000011100110000";
                        f_reg(388) <= "10001111101101010000011011010000";
                        f_reg(389) <= "00010100111101011111111111111100";
                        f_reg(390) <= "10001100000111010000011100110000";
                        f_reg(391) <= "10001111101010000000011011010100";
                        f_reg(392) <= "10001100000111010000011100110000";
                        f_reg(393) <= "10001111101101100000011011010100";
                        f_reg(394) <= "00010101000101101111111111111100";
                        f_reg(395) <= "10001100000111010000011100110000";
                        f_reg(396) <= "10001111101010010000011011011000";
                        f_reg(397) <= "10001100000111010000011100110000";
                        f_reg(398) <= "10001111101101110000011011011000";
                        f_reg(399) <= "00010101001101111111111111111100";
                        f_reg(400) <= "10001100000111010000011100110000";
                        f_reg(401) <= "10001111101010100000011011011100";
                        f_reg(402) <= "10001100000111010000011100110000";
                        f_reg(403) <= "10001111101110000000011011011100";
                        f_reg(404) <= "00010101010110001111111111111100";
                        f_reg(405) <= "10001100000111010000011100110000";
                        f_reg(406) <= "10001111101010110000011011100000";
                        f_reg(407) <= "10001100000111010000011100110000";
                        f_reg(408) <= "10001111101110010000011011100000";
                        f_reg(409) <= "00010101011110011111111111111100";
                        f_reg(410) <= "10001100000111010000011100110000";
                        f_reg(411) <= "10001111101011000000011011100100";
                        f_reg(412) <= "10001100000111010000011100110000";
                        f_reg(413) <= "10001111101110100000011011100100";
                        f_reg(414) <= "00010101100110101111111111111100";
                        f_reg(415) <= "10001100000111010000011100110000";
                        f_reg(416) <= "10001111101011010000011011101000";
                        f_reg(417) <= "10001100000111010000011100110000";
                        f_reg(418) <= "10001111101110110000011011101000";
                        f_reg(419) <= "00010101101110111111111111111100";
                        f_reg(420) <= "10001100000111010000011100110000";
                        f_reg(421) <= "10001111101011100000011011101100";
                        f_reg(422) <= "10001100000111010000011100110000";
                        f_reg(423) <= "10001111101111000000011011101100";
                        f_reg(424) <= "00010101110111001111111111111100";
                        f_reg(425) <= "10001100000111010000011100110000";
                        f_reg(426) <= "10001111101111100000011011110000";
                        f_reg(427) <= "10001100000111010000011100110000";
                        f_reg(428) <= "10001111101111110000011011110000";
                        f_reg(429) <= "00010111110111111111111111111100";
                        f_reg(430) <= "00010000000000001111111100111000";
                        f_reg(431) <= "00000000000000000000000000000000";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000001111100111";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010011010011001001";
                        f_reg(4) <= "00111100000000101001011011000110";
                        f_reg(5) <= "00000000000000010001100000000110";
                        f_reg(6) <= "00101000001001000101110010010011";
                        f_reg(7) <= "10101100000001000000001110101000";
                        f_reg(8) <= "00000000000000000010100000100100";
                        f_reg(9) <= "00000000001000000011000000000110";
                        f_reg(10) <= "00000000110000010011100000100101";
                        f_reg(11) <= "00000000000000000000000000000000";
                        f_reg(12) <= "00000000110000000100000000100010";
                        f_reg(13) <= "00000000000010000100110101000000";
                        f_reg(14) <= "00100100101010101101000010011100";
                        f_reg(15) <= "00000001010001010101100000100011";
                        f_reg(16) <= "00101001011011000011010101010101";
                        f_reg(17) <= "00000000011001000110100000100110";
                        f_reg(18) <= "00000001100001100111000000101010";
                        f_reg(19) <= "00101001110011111011100100100011";
                        f_reg(20) <= "00000000001010111000000000000111";
                        f_reg(21) <= "10101100000010000000001110101100";
                        f_reg(22) <= "00000001101001111000100000000100";
                        f_reg(23) <= "00000000000000000000000000000000";
                        f_reg(24) <= "00000000010000011001000000100101";
                        f_reg(25) <= "00000001011011001001100000100010";
                        f_reg(26) <= "10101100000000100000001110110000";
                        f_reg(27) <= "00000001100011011010000000100101";
                        f_reg(28) <= "00000000000100111010111101000010";
                        f_reg(29) <= "00000010010001111011000000100100";
                        f_reg(30) <= "00110001001101110111010101110011";
                        f_reg(31) <= "00000000000011101100011011000011";
                        f_reg(32) <= "00000000010101011100100000000110";
                        f_reg(33) <= "00000010100001011101000000100011";
                        f_reg(34) <= "00111001110110111101011111110100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000000010100101110000000101010";
                        f_reg(37) <= "10101100000110100000001110110100";
                        f_reg(38) <= "00000010101101101110100000100000";
                        f_reg(39) <= "00000010001010001111000000100110";
                        f_reg(40) <= "00000010000110010101000000100101";
                        f_reg(41) <= "00000011100110000001100000100001";
                        f_reg(42) <= "00000000011010100010000000100000";
                        f_reg(43) <= "00000000000101000011001110000000";
                        f_reg(44) <= "00000010110110000000100000100100";
                        f_reg(45) <= "00000001111111010101100000100110";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00111100000011011000001101011100";
                        f_reg(48) <= "00000010111110011001100000100100";
                        f_reg(49) <= "00000001010110000011100000100010";
                        f_reg(50) <= "00000001100001100100100000000111";
                        f_reg(51) <= "00000001001001000010100000100011";
                        f_reg(52) <= "10101100000110110000001110111000";
                        f_reg(53) <= "00000000111100110111000000100101";
                        f_reg(54) <= "10101100000011100000001110111100";
                        f_reg(55) <= "00000000000001010001000001000000";
                        f_reg(56) <= "00110011110100101010011101011010";
                        f_reg(57) <= "00000001011000101101000000000111";
                        f_reg(58) <= "00000000000000011010110111000000";
                        f_reg(59) <= "00000011101110001000100000101011";
                        f_reg(60) <= "00000010101110100100000000000110";
                        f_reg(61) <= "00100101101100000110000001101101";
                        f_reg(62) <= "00000000000000000000000000000000";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000000000000000000000000000000";
                        f_reg(66) <= "10101100000100000000001111000000";
                        f_reg(67) <= "10101100000100010000001111000100";
                        f_reg(68) <= "10101100000111010000001111001000";
                        f_reg(69) <= "10101100000010000000001111001100";
                        f_reg(70) <= "10101100000100100000001111010000";
                        f_reg(71) <= "00100011111111111111111111111111";
                        f_reg(72) <= "00011111111000001111111110111011";
                        f_reg(73) <= "00010000000000000000000110100111";
                        f_reg(74) <= "00111100000111100000001111100111";
                        f_reg(75) <= "00111100000111110000001111100111";
                        f_reg(76) <= "00000000000111101111010000000010";
                        f_reg(77) <= "00000000000111111111110000000010";
                        f_reg(78) <= "00111100000000010011010011001001";
                        f_reg(79) <= "00111100000011110011010011001001";
                        f_reg(80) <= "00111100000000101001011011000110";
                        f_reg(81) <= "00111100000100001001011011000110";
                        f_reg(82) <= "00000000000000010001100000000110";
                        f_reg(83) <= "00000000000011111000100000000110";
                        f_reg(84) <= "00101000001001000101110010010011";
                        f_reg(85) <= "00101001111100100101110010010011";
                        f_reg(86) <= "00010100100100100000000100001101";
                        f_reg(87) <= "10101100000001000000001110101000";
                        f_reg(88) <= "00000000000000000010100000100100";
                        f_reg(89) <= "00000000000000001001100000100100";
                        f_reg(90) <= "00000000001000000011000000000110";
                        f_reg(91) <= "00000001111000001010000000000110";
                        f_reg(92) <= "00000000110000010011100000100101";
                        f_reg(93) <= "00000010100011111010100000100101";
                        f_reg(94) <= "00000000000000000000000000000000";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000110000000100000000100010";
                        f_reg(97) <= "00000010100000001011000000100010";
                        f_reg(98) <= "00000000000010000100110101000000";
                        f_reg(99) <= "00000000000101101011110101000000";
                        f_reg(100) <= "00100100101010101101000010011100";
                        f_reg(101) <= "00100110011110001101000010011100";
                        f_reg(102) <= "00000001010001010101100000100011";
                        f_reg(103) <= "00000011000100111100100000100011";
                        f_reg(104) <= "00101001011011000011010101010101";
                        f_reg(105) <= "00101011001110100011010101010101";
                        f_reg(106) <= "00000000011001000110100000100110";
                        f_reg(107) <= "00000010001100101101100000100110";
                        f_reg(108) <= "00000001100001100111000000101010";
                        f_reg(109) <= "00000011010101001110000000101010";
                        f_reg(110) <= "00101001110010101011100100100011";
                        f_reg(111) <= "00101011100110001011100100100011";
                        f_reg(112) <= "00000000001010110001100000000111";
                        f_reg(113) <= "00000001111110011000100000000111";
                        f_reg(114) <= "00010101000101100000000011110001";
                        f_reg(115) <= "10101100000010000000001110101100";
                        f_reg(116) <= "00000001101001110010000000000100";
                        f_reg(117) <= "00000011011101011001000000000100";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000010000010011000000100101";
                        f_reg(121) <= "00000010000011111010000000100101";
                        f_reg(122) <= "00000001011011000000100000100010";
                        f_reg(123) <= "00000011001110100111100000100010";
                        f_reg(124) <= "00010100010100000000000011100111";
                        f_reg(125) <= "10101100000000100000001110110000";
                        f_reg(126) <= "00000001100011010101100000100101";
                        f_reg(127) <= "00000011010110111100100000100101";
                        f_reg(128) <= "00000000000000010110111101000010";
                        f_reg(129) <= "00000000000011111101111101000010";
                        f_reg(130) <= "00000000110001110000100000100100";
                        f_reg(131) <= "00000010100101010111100000100100";
                        f_reg(132) <= "00110001001001110111010101110011";
                        f_reg(133) <= "00110010111101010111010101110011";
                        f_reg(134) <= "00000000000011100100111011000011";
                        f_reg(135) <= "00000000000111001011111011000011";
                        f_reg(136) <= "00010101001101110000000011011011";
                        f_reg(137) <= "10101100000010010000001111010100";
                        f_reg(138) <= "00000000010011010100100000000110";
                        f_reg(139) <= "00000010000110111011100000000110";
                        f_reg(140) <= "00010101100110100000000011010111";
                        f_reg(141) <= "10101100000011000000001111011000";
                        f_reg(142) <= "00000001011001010110000000100011";
                        f_reg(143) <= "00000011001100111101000000100011";
                        f_reg(144) <= "00111001110001011101011111110100";
                        f_reg(145) <= "00111011100100111101011111110100";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000010001100111000000101010";
                        f_reg(149) <= "00000010000101001110000000101010";
                        f_reg(150) <= "00010101100110100000000011001101";
                        f_reg(151) <= "10101100000011000000001110110100";
                        f_reg(152) <= "00000001101000010001000000100000";
                        f_reg(153) <= "00000011011011111000000000100000";
                        f_reg(154) <= "00000000100010000011000000100110";
                        f_reg(155) <= "00000010010101101010000000100110";
                        f_reg(156) <= "00000000011010010110000000100101";
                        f_reg(157) <= "00000010001101111101000000100101";
                        f_reg(158) <= "10001100000011010000001111010100";
                        f_reg(159) <= "10001100000110110000001111010100";
                        f_reg(160) <= "00010101101110111111111111111110";
                        f_reg(161) <= "00000001110011010010000000100001";
                        f_reg(162) <= "00000011100110111001000000100001";
                        f_reg(163) <= "00000000100011000100000000100000";
                        f_reg(164) <= "00000010010110101011000000100000";
                        f_reg(165) <= "00000000000010110001101110000000";
                        f_reg(166) <= "00000000000110011000101110000000";
                        f_reg(167) <= "00000000001011010111000000100100";
                        f_reg(168) <= "00000001111110111110000000100100";
                        f_reg(169) <= "00000001010000100010000000100110";
                        f_reg(170) <= "00000011000100001001000000100110";
                        f_reg(171) <= "00000000000000000000000000000000";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00111100000010111000001101011100";
                        f_reg(174) <= "00111100000110011000001101011100";
                        f_reg(175) <= "00000000111010010000100000100100";
                        f_reg(176) <= "00000010101101110111100000100100";
                        f_reg(177) <= "00000001100011010101000000100010";
                        f_reg(178) <= "00000011010110111100000000100010";
                        f_reg(179) <= "10001100000001110000001111011000";
                        f_reg(180) <= "10001100000101010000001111011000";
                        f_reg(181) <= "00010100111101011111111111111110";
                        f_reg(182) <= "00000000111000110100100000000111";
                        f_reg(183) <= "00000010101100011011100000000111";
                        f_reg(184) <= "00000001001010000110000000100011";
                        f_reg(185) <= "00000010111101101101000000100011";
                        f_reg(186) <= "00010100101100110000000010101001";
                        f_reg(187) <= "10101100000001010000001110111000";
                        f_reg(188) <= "00000001010000010001100000100101";
                        f_reg(189) <= "00000011000011111000100000100101";
                        f_reg(190) <= "00010100011100010000000010100101";
                        f_reg(191) <= "10101100000000110000001110111100";
                        f_reg(192) <= "00000000000011000011100001000000";
                        f_reg(193) <= "00000000000110101010100001000000";
                        f_reg(194) <= "00110000110010011010011101011010";
                        f_reg(195) <= "00110010100101111010011101011010";
                        f_reg(196) <= "00000000100001110100000000000111";
                        f_reg(197) <= "00000010010101011011000000000111";
                        f_reg(198) <= "00000000000011100010110111000000";
                        f_reg(199) <= "00000000000111001001110111000000";
                        f_reg(200) <= "00000000010011010101000000101011";
                        f_reg(201) <= "00000010000110111100000000101011";
                        f_reg(202) <= "00000000101010000000100000000110";
                        f_reg(203) <= "00000010011101100111100000000110";
                        f_reg(204) <= "00100101011000110110000001101101";
                        f_reg(205) <= "00100111001100010110000001101101";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00010100011100010000000010001101";
                        f_reg(215) <= "10101100000000110000001111000000";
                        f_reg(216) <= "00010101010110000000000010001011";
                        f_reg(217) <= "10101100000010100000001111000100";
                        f_reg(218) <= "00010100010100000000000010001001";
                        f_reg(219) <= "10101100000000100000001111001000";
                        f_reg(220) <= "00010100001011110000000010000111";
                        f_reg(221) <= "10101100000000010000001111001100";
                        f_reg(222) <= "00010101001101110000000010000101";
                        f_reg(223) <= "10101100000010010000001111010000";
                        f_reg(224) <= "00100011110111011111111100000110";
                        f_reg(225) <= "00010011101000000000000000010111";
                        f_reg(226) <= "00100011110111011111111000001100";
                        f_reg(227) <= "00010011101000000000000000010101";
                        f_reg(228) <= "00100011110111011111110100010010";
                        f_reg(229) <= "00010011101000000000000000010011";
                        f_reg(230) <= "00100011110111101111111111111111";
                        f_reg(231) <= "00100011111111111111111111111111";
                        f_reg(232) <= "00010111110111110000000001111011";
                        f_reg(233) <= "00011111111000001111111101100101";
                        f_reg(234) <= "00010000000000000000000100000110";
                        f_reg(235) <= "00000000000000000000000000000000";
                        f_reg(236) <= "00000000000000000000000000000000";
                        f_reg(237) <= "00000000000000000000000000000000";
                        f_reg(238) <= "00000000000000000000000000000000";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000000000000000000000000000000";
                        f_reg(242) <= "00000000000000000000000000000000";
                        f_reg(243) <= "00000000000000000000000000000000";
                        f_reg(244) <= "00000000000000000000000000000000";
                        f_reg(245) <= "00000000000000000000000000000000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "10001100000111010000011100110000";
                        f_reg(249) <= "00011111101000000000000000000011";
                        f_reg(250) <= "00100000000111010000000000111100";
                        f_reg(251) <= "00010000000000000000000000000010";
                        f_reg(252) <= "00100000000111010000000000000000";
                        f_reg(253) <= "00010100001011110000000001100110";
                        f_reg(254) <= "10101111101000010000011010111000";
                        f_reg(255) <= "10001100000111010000011100110000";
                        f_reg(256) <= "00011111101000000000000000000011";
                        f_reg(257) <= "00100000000111010000000000111100";
                        f_reg(258) <= "00010000000000000000000000000010";
                        f_reg(259) <= "00100000000111010000000000000000";
                        f_reg(260) <= "00010100010100000000000001011111";
                        f_reg(261) <= "10101111101000100000011010111100";
                        f_reg(262) <= "10001100000111010000011100110000";
                        f_reg(263) <= "00011111101000000000000000000011";
                        f_reg(264) <= "00100000000111010000000000111100";
                        f_reg(265) <= "00010000000000000000000000000010";
                        f_reg(266) <= "00100000000111010000000000000000";
                        f_reg(267) <= "00010100011100010000000001011000";
                        f_reg(268) <= "10101111101000110000011011000000";
                        f_reg(269) <= "10001100000111010000011100110000";
                        f_reg(270) <= "00011111101000000000000000000011";
                        f_reg(271) <= "00100000000111010000000000111100";
                        f_reg(272) <= "00010000000000000000000000000010";
                        f_reg(273) <= "00100000000111010000000000000000";
                        f_reg(274) <= "00010100100100100000000001010001";
                        f_reg(275) <= "10101111101001000000011011000100";
                        f_reg(276) <= "10001100000111010000011100110000";
                        f_reg(277) <= "00011111101000000000000000000011";
                        f_reg(278) <= "00100000000111010000000000111100";
                        f_reg(279) <= "00010000000000000000000000000010";
                        f_reg(280) <= "00100000000111010000000000000000";
                        f_reg(281) <= "00010100101100110000000001001010";
                        f_reg(282) <= "10101111101001010000011011001000";
                        f_reg(283) <= "10001100000111010000011100110000";
                        f_reg(284) <= "00011111101000000000000000000011";
                        f_reg(285) <= "00100000000111010000000000111100";
                        f_reg(286) <= "00010000000000000000000000000010";
                        f_reg(287) <= "00100000000111010000000000000000";
                        f_reg(288) <= "00010100110101000000000001000011";
                        f_reg(289) <= "10101111101001100000011011001100";
                        f_reg(290) <= "10001100000111010000011100110000";
                        f_reg(291) <= "00011111101000000000000000000011";
                        f_reg(292) <= "00100000000111010000000000111100";
                        f_reg(293) <= "00010000000000000000000000000010";
                        f_reg(294) <= "00100000000111010000000000000000";
                        f_reg(295) <= "00010100111101010000000000111100";
                        f_reg(296) <= "10101111101001110000011011010000";
                        f_reg(297) <= "10001100000111010000011100110000";
                        f_reg(298) <= "00011111101000000000000000000011";
                        f_reg(299) <= "00100000000111010000000000111100";
                        f_reg(300) <= "00010000000000000000000000000010";
                        f_reg(301) <= "00100000000111010000000000000000";
                        f_reg(302) <= "00010101000101100000000000110101";
                        f_reg(303) <= "10101111101010000000011011010100";
                        f_reg(304) <= "10001100000111010000011100110000";
                        f_reg(305) <= "00011111101000000000000000000011";
                        f_reg(306) <= "00100000000111010000000000111100";
                        f_reg(307) <= "00010000000000000000000000000010";
                        f_reg(308) <= "00100000000111010000000000000000";
                        f_reg(309) <= "00010101001101110000000000101110";
                        f_reg(310) <= "10101111101010010000011011011000";
                        f_reg(311) <= "10001100000111010000011100110000";
                        f_reg(312) <= "00011111101000000000000000000011";
                        f_reg(313) <= "00100000000111010000000000111100";
                        f_reg(314) <= "00010000000000000000000000000010";
                        f_reg(315) <= "00100000000111010000000000000000";
                        f_reg(316) <= "00010101010110000000000000100111";
                        f_reg(317) <= "10101111101010100000011011011100";
                        f_reg(318) <= "10001100000111010000011100110000";
                        f_reg(319) <= "00011111101000000000000000000011";
                        f_reg(320) <= "00100000000111010000000000111100";
                        f_reg(321) <= "00010000000000000000000000000010";
                        f_reg(322) <= "00100000000111010000000000000000";
                        f_reg(323) <= "00010101011110010000000000100000";
                        f_reg(324) <= "10101111101010110000011011100000";
                        f_reg(325) <= "10001100000111010000011100110000";
                        f_reg(326) <= "00011111101000000000000000000011";
                        f_reg(327) <= "00100000000111010000000000111100";
                        f_reg(328) <= "00010000000000000000000000000010";
                        f_reg(329) <= "00100000000111010000000000000000";
                        f_reg(330) <= "00010101100110100000000000011001";
                        f_reg(331) <= "10101111101011000000011011100100";
                        f_reg(332) <= "10001100000111010000011100110000";
                        f_reg(333) <= "00011111101000000000000000000011";
                        f_reg(334) <= "00100000000111010000000000111100";
                        f_reg(335) <= "00010000000000000000000000000010";
                        f_reg(336) <= "00100000000111010000000000000000";
                        f_reg(337) <= "00010101101110110000000000010010";
                        f_reg(338) <= "10101111101011010000011011101000";
                        f_reg(339) <= "10001100000111010000011100110000";
                        f_reg(340) <= "00011111101000000000000000000011";
                        f_reg(341) <= "00100000000111010000000000111100";
                        f_reg(342) <= "00010000000000000000000000000010";
                        f_reg(343) <= "00100000000111010000000000000000";
                        f_reg(344) <= "00010101110111000000000000001011";
                        f_reg(345) <= "10101111101011100000011011101100";
                        f_reg(346) <= "10001100000111010000011100110000";
                        f_reg(347) <= "00011111101000000000000000000011";
                        f_reg(348) <= "00100000000111010000000000111100";
                        f_reg(349) <= "00010000000000000000000000000010";
                        f_reg(350) <= "00100000000111010000000000000000";
                        f_reg(351) <= "00010111110111110000000000000100";
                        f_reg(352) <= "10101111101111100000011011110000";
                        f_reg(353) <= "10101100000111010000011100110000";
                        f_reg(354) <= "00010000000000001111111110000100";
                        f_reg(355) <= "10001100000111010000011100110000";
                        f_reg(356) <= "10001111101000010000011010111000";
                        f_reg(357) <= "10001100000111010000011100110000";
                        f_reg(358) <= "10001111101011110000011010111000";
                        f_reg(359) <= "00010100001011111111111111111100";
                        f_reg(360) <= "10001100000111010000011100110000";
                        f_reg(361) <= "10001111101000100000011010111100";
                        f_reg(362) <= "10001100000111010000011100110000";
                        f_reg(363) <= "10001111101100000000011010111100";
                        f_reg(364) <= "00010100010100001111111111111100";
                        f_reg(365) <= "10001100000111010000011100110000";
                        f_reg(366) <= "10001111101000110000011011000000";
                        f_reg(367) <= "10001100000111010000011100110000";
                        f_reg(368) <= "10001111101100010000011011000000";
                        f_reg(369) <= "00010100011100011111111111111100";
                        f_reg(370) <= "10001100000111010000011100110000";
                        f_reg(371) <= "10001111101001000000011011000100";
                        f_reg(372) <= "10001100000111010000011100110000";
                        f_reg(373) <= "10001111101100100000011011000100";
                        f_reg(374) <= "00010100100100101111111111111100";
                        f_reg(375) <= "10001100000111010000011100110000";
                        f_reg(376) <= "10001111101001010000011011001000";
                        f_reg(377) <= "10001100000111010000011100110000";
                        f_reg(378) <= "10001111101100110000011011001000";
                        f_reg(379) <= "00010100101100111111111111111100";
                        f_reg(380) <= "10001100000111010000011100110000";
                        f_reg(381) <= "10001111101001100000011011001100";
                        f_reg(382) <= "10001100000111010000011100110000";
                        f_reg(383) <= "10001111101101000000011011001100";
                        f_reg(384) <= "00010100110101001111111111111100";
                        f_reg(385) <= "10001100000111010000011100110000";
                        f_reg(386) <= "10001111101001110000011011010000";
                        f_reg(387) <= "10001100000111010000011100110000";
                        f_reg(388) <= "10001111101101010000011011010000";
                        f_reg(389) <= "00010100111101011111111111111100";
                        f_reg(390) <= "10001100000111010000011100110000";
                        f_reg(391) <= "10001111101010000000011011010100";
                        f_reg(392) <= "10001100000111010000011100110000";
                        f_reg(393) <= "10001111101101100000011011010100";
                        f_reg(394) <= "00010101000101101111111111111100";
                        f_reg(395) <= "10001100000111010000011100110000";
                        f_reg(396) <= "10001111101010010000011011011000";
                        f_reg(397) <= "10001100000111010000011100110000";
                        f_reg(398) <= "10001111101101110000011011011000";
                        f_reg(399) <= "00010101001101111111111111111100";
                        f_reg(400) <= "10001100000111010000011100110000";
                        f_reg(401) <= "10001111101010100000011011011100";
                        f_reg(402) <= "10001100000111010000011100110000";
                        f_reg(403) <= "10001111101110000000011011011100";
                        f_reg(404) <= "00010101010110001111111111111100";
                        f_reg(405) <= "10001100000111010000011100110000";
                        f_reg(406) <= "10001111101010110000011011100000";
                        f_reg(407) <= "10001100000111010000011100110000";
                        f_reg(408) <= "10001111101110010000011011100000";
                        f_reg(409) <= "00010101011110011111111111111100";
                        f_reg(410) <= "10001100000111010000011100110000";
                        f_reg(411) <= "10001111101011000000011011100100";
                        f_reg(412) <= "10001100000111010000011100110000";
                        f_reg(413) <= "10001111101110100000011011100100";
                        f_reg(414) <= "00010101100110101111111111111100";
                        f_reg(415) <= "10001100000111010000011100110000";
                        f_reg(416) <= "10001111101011010000011011101000";
                        f_reg(417) <= "10001100000111010000011100110000";
                        f_reg(418) <= "10001111101110110000011011101000";
                        f_reg(419) <= "00010101101110111111111111111100";
                        f_reg(420) <= "10001100000111010000011100110000";
                        f_reg(421) <= "10001111101011100000011011101100";
                        f_reg(422) <= "10001100000111010000011100110000";
                        f_reg(423) <= "10001111101111000000011011101100";
                        f_reg(424) <= "00010101110111001111111111111100";
                        f_reg(425) <= "10001100000111010000011100110000";
                        f_reg(426) <= "10001111101111100000011011110000";
                        f_reg(427) <= "10001100000111010000011100110000";
                        f_reg(428) <= "10001111101111110000011011110000";
                        f_reg(429) <= "00010111110111111111111111111100";
                        f_reg(430) <= "00010000000000001111111100111000";
                        f_reg(431) <= "00000000000000000000000000000000";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000001111100111";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 13513
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- LUI R2 -26938
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SRLV R3 R1 R0
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SLTI R4 R1 23699
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SW R4 R0 936
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- AND R5 R0 R0
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- SRLV R6 R0 R1
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- OR R7 R6 R1
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- NOP
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- SUB R8 R6 R0
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- SLL R9 R8 21
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- ADDIU R10 R5 -12132
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- SUBU R11 R10 R5
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- SLTI R12 R11 13653
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- XOR R13 R3 R4
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- SLT R14 R12 R6
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SLTI R15 R14 -18141
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- SRAV R16 R11 R1
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SW R8 R0 940
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- SLLV R17 R7 R13
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- NOP
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- OR R18 R2 R1
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- SUB R19 R11 R12
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- SW R2 R0 944
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- OR R20 R12 R13
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- SRL R21 R19 29
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- AND R22 R18 R7
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- ANDI R23 R9 30067
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- SRA R24 R14 27
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- SRLV R25 R21 R2
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- SUBU R26 R20 R5
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- XORI R27 R14 -10252
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- NOP
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- SLT R28 R2 R18
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- SW R26 R0 948
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- ADD R29 R21 R22
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- XOR R30 R17 R8
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- OR R10 R16 R25
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- ADDU R3 R28 R24
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- ADD R4 R3 R10
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SLL R6 R20 14
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- AND R1 R22 R24
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- XOR R11 R15 R29
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- NOP
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- LUI R13 -31908
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- AND R19 R23 R25
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- SUB R7 R10 R24
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- SRAV R9 R6 R12
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SUBU R5 R9 R4
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- SW R27 R0 952
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- OR R14 R7 R19
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SW R14 R0 956
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SLL R2 R5 1
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- ANDI R18 R30 -22694
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SRAV R26 R2 R11
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- SLL R21 R1 23
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- SLTU R17 R29 R24
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SRLV R8 R26 R21
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- ADDIU R16 R13 24685
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- NOP
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- NOP
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- NOP
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- NOP
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- SW R16 R0 960
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- SW R17 R0 964
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- SW R29 R0 968
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- SW R8 R0 972
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SW R18 R0 976
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- ADDI R31 R31 -1
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- BGTZ R31 -69
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- BEQ R0 R0 423
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- LUI R30 999
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- LUI R31 999
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- SRL R30 R30 16
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- SRL R31 R31 16
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- LUI R1 13513
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- LUI R15 13513
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- LUI R2 -26938
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- LUI R16 -26938
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- SRLV R3 R1 R0
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SRLV R17 R15 R0
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- SLTI R4 R1 23699
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- SLTI R18 R15 23699
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- BNE R4 R18 269
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SW R4 R0 936
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- AND R5 R0 R0
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- AND R19 R0 R0
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- SRLV R6 R0 R1
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- SRLV R20 R0 R15
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- OR R7 R6 R1
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- OR R21 R20 R15
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- NOP
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- NOP
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- SUB R8 R6 R0
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SUB R22 R20 R0
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SLL R9 R8 21
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- SLL R23 R22 21
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- ADDIU R10 R5 -12132
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- ADDIU R24 R19 -12132
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- SUBU R11 R10 R5
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SUBU R25 R24 R19
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- SLTI R12 R11 13653
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- SLTI R26 R25 13653
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- XOR R13 R3 R4
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- XOR R27 R17 R18
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- SLT R14 R12 R6
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- SLT R28 R26 R20
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- SLTI R10 R14 -18141
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- SLTI R24 R28 -18141
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- SRAV R3 R11 R1
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- SRAV R17 R25 R15
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- BNE R8 R22 241
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- SW R8 R0 940
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- SLLV R4 R7 R13
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- SLLV R18 R21 R27
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- NOP
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- NOP
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- OR R6 R2 R1
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- OR R20 R16 R15
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- SUB R1 R11 R12
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- SUB R15 R25 R26
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- BNE R2 R16 231
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- SW R2 R0 944
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- OR R11 R12 R13
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- OR R25 R26 R27
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SRL R13 R1 29
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- SRL R27 R15 29
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- AND R1 R6 R7
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- AND R15 R20 R21
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- ANDI R7 R9 30067
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- ANDI R21 R23 30067
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- SRA R9 R14 27
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- SRA R23 R28 27
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- BNE R9 R23 219
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- SW R9 R0 980
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SRLV R9 R13 R2
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- SRLV R23 R27 R16
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- BNE R12 R26 215
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- SW R12 R0 984
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- SUBU R12 R11 R5
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- SUBU R26 R25 R19
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- XORI R5 R14 -10252
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- XORI R19 R28 -10252
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- NOP
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- NOP
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- SLT R14 R2 R6
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- SLT R28 R16 R20
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- BNE R12 R26 205
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- SW R12 R0 948
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- ADD R2 R13 R1
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- ADD R16 R27 R15
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- XOR R6 R4 R8
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- XOR R20 R18 R22
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- OR R12 R3 R9
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- OR R26 R17 R23
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- LW R13 R0 980
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- LW R27 R0 980
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- BNE R13 R27 -2
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- ADDU R4 R14 R13
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- ADDU R18 R28 R27
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- ADD R8 R4 R12
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- ADD R22 R18 R26
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- SLL R3 R11 14
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- SLL R17 R25 14
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- AND R14 R1 R13
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- AND R28 R15 R27
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- XOR R4 R10 R2
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- XOR R18 R24 R16
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- NOP
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- NOP
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- LUI R11 -31908
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- LUI R25 -31908
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- AND R1 R7 R9
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- AND R15 R21 R23
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- SUB R10 R12 R13
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- SUB R24 R26 R27
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- LW R7 R0 984
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- LW R21 R0 984
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- BNE R7 R21 -2
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SRAV R9 R3 R7
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- SRAV R23 R17 R21
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- SUBU R12 R9 R8
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- SUBU R26 R23 R22
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- BNE R5 R19 169
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- SW R5 R0 952
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- OR R3 R10 R1
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- OR R17 R24 R15
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- BNE R3 R17 165
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- SW R3 R0 956
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- SLL R7 R12 1
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- SLL R21 R26 1
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- ANDI R9 R6 -22694
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- ANDI R23 R20 -22694
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- SRAV R8 R7 R4
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- SRAV R22 R21 R18
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- SLL R5 R14 23
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- SLL R19 R28 23
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- SLTU R10 R2 R13
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- SLTU R24 R16 R27
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- SRLV R1 R8 R5
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- SRLV R15 R22 R19
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- ADDIU R3 R11 24685
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- ADDIU R17 R25 24685
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- NOP
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- NOP
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- NOP
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- NOP
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- NOP
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- NOP
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- NOP
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- NOP
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- BNE R3 R17 141
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- SW R3 R0 960
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- BNE R10 R24 139
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- SW R10 R0 964
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- BNE R2 R16 137
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- SW R2 R0 968
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- BNE R1 R15 135
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- SW R1 R0 972
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- BNE R9 R23 133
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- SW R9 R0 976
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- ADDI R29 R30 -250
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- BEQ R29 R0 23
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- ADDI R29 R30 -500
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- BEQ R29 R0 21
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- ADDI R29 R30 -750
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- BEQ R29 R0 19
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- ADDI R30 R30 -1
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- ADDI R31 R31 -1
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- BNE R30 R31 123
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- BGTZ R31 -155
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- BEQ R0 R0 262
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- NOP
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- NOP
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- NOP
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- NOP
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- NOP
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- NOP
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- NOP
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- NOP
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- NOP
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- NOP
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- NOP
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- NOP
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- NOP
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- LW R29 R0 1840
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- BGTZ R29 3
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- ADDI R29 R0 60
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- BEQ R0 R0 2
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- ADDI R29 R0 0
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- BNE R1 R15 102
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- SW R1 R29 1720
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- LW R29 R0 1840
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- BGTZ R29 3
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- ADDI R29 R0 60
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- BEQ R0 R0 2
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- ADDI R29 R0 0
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- BNE R2 R16 95
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- SW R2 R29 1724
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- LW R29 R0 1840
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- BGTZ R29 3
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- ADDI R29 R0 60
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- BEQ R0 R0 2
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- ADDI R29 R0 0
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- BNE R3 R17 88
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- SW R3 R29 1728
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- LW R29 R0 1840
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- BGTZ R29 3
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- ADDI R29 R0 60
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- BEQ R0 R0 2
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- ADDI R29 R0 0
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- BNE R4 R18 81
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- SW R4 R29 1732
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- LW R29 R0 1840
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- BGTZ R29 3
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- ADDI R29 R0 60
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- BEQ R0 R0 2
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- ADDI R29 R0 0
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- BNE R5 R19 74
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- SW R5 R29 1736
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- LW R29 R0 1840
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- BGTZ R29 3
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- ADDI R29 R0 60
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- BEQ R0 R0 2
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- ADDI R29 R0 0
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- BNE R6 R20 67
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- SW R6 R29 1740
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- LW R29 R0 1840
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- BGTZ R29 3
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- ADDI R29 R0 60
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- BEQ R0 R0 2
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- ADDI R29 R0 0
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- BNE R7 R21 60
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- SW R7 R29 1744
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- LW R29 R0 1840
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- BGTZ R29 3
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- ADDI R29 R0 60
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- BEQ R0 R0 2
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- ADDI R29 R0 0
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- BNE R8 R22 53
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- SW R8 R29 1748
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- LW R29 R0 1840
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- BGTZ R29 3
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- ADDI R29 R0 60
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- BEQ R0 R0 2
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- ADDI R29 R0 0
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- BNE R9 R23 46
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- SW R9 R29 1752
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- LW R29 R0 1840
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- BGTZ R29 3
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- ADDI R29 R0 60
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- BEQ R0 R0 2
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- ADDI R29 R0 0
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- BNE R10 R24 39
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- SW R10 R29 1756
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- LW R29 R0 1840
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- BGTZ R29 3
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- ADDI R29 R0 60
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- BEQ R0 R0 2
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- ADDI R29 R0 0
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- BNE R11 R25 32
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- SW R11 R29 1760
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- LW R29 R0 1840
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- BGTZ R29 3
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- ADDI R29 R0 60
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- BEQ R0 R0 2
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- ADDI R29 R0 0
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- BNE R12 R26 25
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- SW R12 R29 1764
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- LW R29 R0 1840
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- BGTZ R29 3
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- ADDI R29 R0 60
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- BEQ R0 R0 2
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- ADDI R29 R0 0
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- BNE R13 R27 18
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- SW R13 R29 1768
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- LW R29 R0 1840
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- BGTZ R29 3
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- ADDI R29 R0 60
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- BEQ R0 R0 2
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- ADDI R29 R0 0
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- BNE R14 R28 11
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- SW R14 R29 1772
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- LW R29 R0 1840
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- BGTZ R29 3
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- ADDI R29 R0 60
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- BEQ R0 R0 2
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- ADDI R29 R0 0
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- BNE R30 R31 4
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- SW R30 R29 1776
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- SW R29 R0 1840
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- BEQ R0 R0 -124
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- LW R29 R0 1840
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- LW R1 R29 1720
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- LW R29 R0 1840
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- LW R15 R29 1720
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- BNE R1 R15 -4
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- LW R29 R0 1840
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- LW R2 R29 1724
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- LW R29 R0 1840
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- LW R16 R29 1724
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- BNE R2 R16 -4
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- LW R29 R0 1840
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- LW R3 R29 1728
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- LW R29 R0 1840
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- LW R17 R29 1728
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- BNE R3 R17 -4
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- LW R29 R0 1840
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- LW R4 R29 1732
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- LW R29 R0 1840
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- LW R18 R29 1732
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- BNE R4 R18 -4
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- LW R29 R0 1840
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- LW R5 R29 1736
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- LW R29 R0 1840
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- LW R19 R29 1736
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- BNE R5 R19 -4
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- LW R29 R0 1840
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- LW R6 R29 1740
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- LW R29 R0 1840
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- LW R20 R29 1740
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- BNE R6 R20 -4
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- LW R29 R0 1840
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- LW R7 R29 1744
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- LW R29 R0 1840
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- LW R21 R29 1744
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- BNE R7 R21 -4
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- LW R29 R0 1840
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- LW R8 R29 1748
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- LW R29 R0 1840
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- LW R22 R29 1748
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- BNE R8 R22 -4
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- LW R29 R0 1840
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- LW R9 R29 1752
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- LW R29 R0 1840
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- LW R23 R29 1752
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- BNE R9 R23 -4
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- LW R29 R0 1840
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- LW R10 R29 1756
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- LW R29 R0 1840
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- LW R24 R29 1756
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- BNE R10 R24 -4
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- LW R29 R0 1840
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- LW R11 R29 1760
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- LW R29 R0 1840
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- LW R25 R29 1760
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- BNE R11 R25 -4
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- LW R29 R0 1840
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- LW R12 R29 1764
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- LW R29 R0 1840
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- LW R26 R29 1764
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- BNE R12 R26 -4
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- LW R29 R0 1840
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- LW R13 R29 1768
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- LW R29 R0 1840
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- LW R27 R29 1768
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- BNE R13 R27 -4
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- LW R29 R0 1840
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- LW R14 R29 1772
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- LW R29 R0 1840
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- LW R28 R29 1772
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- BNE R14 R28 -4
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R29 R0 1840
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R30 R29 1776
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- LW R29 R0 1840
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- LW R31 R29 1776
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- BNE R30 R31 -4
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- BEQ R0 R0 -200
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- NOP
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- NOP
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- NOP
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- NOP
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- NOP
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- NOP
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- NOP
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- NOP
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- NOP
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- NOP
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- NOP
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- NOP
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- NOP
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- NOP
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- NOP
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- NOP
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- NOP
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- NOP
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- NOP
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- NOP
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- NOP
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- NOP
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- NOP
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- NOP
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- NOP
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- NOP
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- NOP
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- NOP
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- NOP
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- NOP
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- NOP
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- NOP
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- NOP
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- NOP
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- NOP
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- NOP
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- NOP
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- NOP
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- NOP
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- NOP
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- NOP
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- NOP
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- NOP
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- NOP
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- NOP
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- NOP
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- NOP
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- NOP
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- NOP
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- NOP
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- NOP
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- NOP
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- NOP
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- NOP
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- NOP
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- NOP
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- NOP
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- NOP
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- NOP
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- NOP
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- NOP
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- NOP
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- NOP
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- NOP
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- NOP
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010011010011001001";
                        f_reg(4) <= "00111100000000101001011011000110";
                        f_reg(5) <= "00000000000000010001100000000110";
                        f_reg(6) <= "00101000001001000101110010010011";
                        f_reg(7) <= "10101100000001000000001110101000";
                        f_reg(8) <= "00000000000000000010100000100100";
                        f_reg(9) <= "00000000001000000011000000000110";
                        f_reg(10) <= "00000000110000010011100000100101";
                        f_reg(11) <= "00000000000000000000000000000000";
                        f_reg(12) <= "00000000110000000100000000100010";
                        f_reg(13) <= "00000000000010000100110101000000";
                        f_reg(14) <= "00100100101010101101000010011100";
                        f_reg(15) <= "00000001010001010101100000100011";
                        f_reg(16) <= "00101001011011000011010101010101";
                        f_reg(17) <= "00000000011001000110100000100110";
                        f_reg(18) <= "00000001100001100111000000101010";
                        f_reg(19) <= "00101001110011111011100100100011";
                        f_reg(20) <= "00000000001010111000000000000111";
                        f_reg(21) <= "10101100000010000000001110101100";
                        f_reg(22) <= "00000001101001111000100000000100";
                        f_reg(23) <= "00000000000000000000000000000000";
                        f_reg(24) <= "00000000010000011001000000100101";
                        f_reg(25) <= "00000001011011001001100000100010";
                        f_reg(26) <= "10101100000000100000001110110000";
                        f_reg(27) <= "00000001100011011010000000100101";
                        f_reg(28) <= "00000000000100111010111101000010";
                        f_reg(29) <= "00000010010001111011000000100100";
                        f_reg(30) <= "00110001001101110111010101110011";
                        f_reg(31) <= "00000000000011101100011011000011";
                        f_reg(32) <= "00000000010101011100100000000110";
                        f_reg(33) <= "00000010100001011101000000100011";
                        f_reg(34) <= "00111001110110111101011111110100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000000010100101110000000101010";
                        f_reg(37) <= "10101100000110100000001110110100";
                        f_reg(38) <= "00000010101101101110100000100000";
                        f_reg(39) <= "00000010001010001111000000100110";
                        f_reg(40) <= "00000010000110010101000000100101";
                        f_reg(41) <= "00000011100110000001100000100001";
                        f_reg(42) <= "00000000011010100010000000100000";
                        f_reg(43) <= "00000000000101000011001110000000";
                        f_reg(44) <= "00000010110110000000100000100100";
                        f_reg(45) <= "00000001111111010101100000100110";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00111100000011011000001101011100";
                        f_reg(48) <= "00000010111110011001100000100100";
                        f_reg(49) <= "00000001010110000011100000100010";
                        f_reg(50) <= "00000001100001100100100000000111";
                        f_reg(51) <= "00000001001001000010100000100011";
                        f_reg(52) <= "10101100000110110000001110111000";
                        f_reg(53) <= "00000000111100110111000000100101";
                        f_reg(54) <= "10101100000011100000001110111100";
                        f_reg(55) <= "00000000000001010001000001000000";
                        f_reg(56) <= "00110011110100101010011101011010";
                        f_reg(57) <= "00000001011000101101000000000111";
                        f_reg(58) <= "00000000000000011010110111000000";
                        f_reg(59) <= "00000011101110001000100000101011";
                        f_reg(60) <= "00000010101110100100000000000110";
                        f_reg(61) <= "00100101101100000110000001101101";
                        f_reg(62) <= "00000000000000000000000000000000";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000000000000000000000000000000";
                        f_reg(66) <= "10101100000100000000001111000000";
                        f_reg(67) <= "10101100000100010000001111000100";
                        f_reg(68) <= "10101100000111010000001111001000";
                        f_reg(69) <= "10101100000010000000001111001100";
                        f_reg(70) <= "10101100000100100000001111010000";
                        f_reg(71) <= "00100011111111111111111111111111";
                        f_reg(72) <= "00011111111000001111111110111011";
                        f_reg(73) <= "00010000000000000000000110100111";
                        f_reg(74) <= "00111100000111100000001111100111";
                        f_reg(75) <= "00111100000111110000001111100111";
                        f_reg(76) <= "00000000000111101111010000000010";
                        f_reg(77) <= "00000000000111111111110000000010";
                        f_reg(78) <= "00111100000000010011010011001001";
                        f_reg(79) <= "00111100000011110011010011001001";
                        f_reg(80) <= "00111100000000101001011011000110";
                        f_reg(81) <= "00111100000100001001011011000110";
                        f_reg(82) <= "00000000000000010001100000000110";
                        f_reg(83) <= "00000000000011111000100000000110";
                        f_reg(84) <= "00101000001001000101110010010011";
                        f_reg(85) <= "00101001111100100101110010010011";
                        f_reg(86) <= "00010100100100100000000100001101";
                        f_reg(87) <= "10101100000001000000001110101000";
                        f_reg(88) <= "00000000000000000010100000100100";
                        f_reg(89) <= "00000000000000001001100000100100";
                        f_reg(90) <= "00000000001000000011000000000110";
                        f_reg(91) <= "00000001111000001010000000000110";
                        f_reg(92) <= "00000000110000010011100000100101";
                        f_reg(93) <= "00000010100011111010100000100101";
                        f_reg(94) <= "00000000000000000000000000000000";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000110000000100000000100010";
                        f_reg(97) <= "00000010100000001011000000100010";
                        f_reg(98) <= "00000000000010000100110101000000";
                        f_reg(99) <= "00000000000101101011110101000000";
                        f_reg(100) <= "00100100101010101101000010011100";
                        f_reg(101) <= "00100110011110001101000010011100";
                        f_reg(102) <= "00000001010001010101100000100011";
                        f_reg(103) <= "00000011000100111100100000100011";
                        f_reg(104) <= "00101001011011000011010101010101";
                        f_reg(105) <= "00101011001110100011010101010101";
                        f_reg(106) <= "00000000011001000110100000100110";
                        f_reg(107) <= "00000010001100101101100000100110";
                        f_reg(108) <= "00000001100001100111000000101010";
                        f_reg(109) <= "00000011010101001110000000101010";
                        f_reg(110) <= "00101001110010101011100100100011";
                        f_reg(111) <= "00101011100110001011100100100011";
                        f_reg(112) <= "00000000001010110001100000000111";
                        f_reg(113) <= "00000001111110011000100000000111";
                        f_reg(114) <= "00010101000101100000000011110001";
                        f_reg(115) <= "10101100000010000000001110101100";
                        f_reg(116) <= "00000001101001110010000000000100";
                        f_reg(117) <= "00000011011101011001000000000100";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000010000010011000000100101";
                        f_reg(121) <= "00000010000011111010000000100101";
                        f_reg(122) <= "00000001011011000000100000100010";
                        f_reg(123) <= "00000011001110100111100000100010";
                        f_reg(124) <= "00010100010100000000000011100111";
                        f_reg(125) <= "10101100000000100000001110110000";
                        f_reg(126) <= "00000001100011010101100000100101";
                        f_reg(127) <= "00000011010110111100100000100101";
                        f_reg(128) <= "00000000000000010110111101000010";
                        f_reg(129) <= "00000000000011111101111101000010";
                        f_reg(130) <= "00000000110001110000100000100100";
                        f_reg(131) <= "00000010100101010111100000100100";
                        f_reg(132) <= "00110001001001110111010101110011";
                        f_reg(133) <= "00110010111101010111010101110011";
                        f_reg(134) <= "00000000000011100100111011000011";
                        f_reg(135) <= "00000000000111001011111011000011";
                        f_reg(136) <= "00010101001101110000000011011011";
                        f_reg(137) <= "10101100000010010000001111010100";
                        f_reg(138) <= "00000000010011010100100000000110";
                        f_reg(139) <= "00000010000110111011100000000110";
                        f_reg(140) <= "00010101100110100000000011010111";
                        f_reg(141) <= "10101100000011000000001111011000";
                        f_reg(142) <= "00000001011001010110000000100011";
                        f_reg(143) <= "00000011001100111101000000100011";
                        f_reg(144) <= "00111001110001011101011111110100";
                        f_reg(145) <= "00111011100100111101011111110100";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000010001100111000000101010";
                        f_reg(149) <= "00000010000101001110000000101010";
                        f_reg(150) <= "00010101100110100000000011001101";
                        f_reg(151) <= "10101100000011000000001110110100";
                        f_reg(152) <= "00000001101000010001000000100000";
                        f_reg(153) <= "00000011011011111000000000100000";
                        f_reg(154) <= "00000000100010000011000000100110";
                        f_reg(155) <= "00000010010101101010000000100110";
                        f_reg(156) <= "00000000011010010110000000100101";
                        f_reg(157) <= "00000010001101111101000000100101";
                        f_reg(158) <= "10001100000011010000001111010100";
                        f_reg(159) <= "10001100000110110000001111010100";
                        f_reg(160) <= "00010101101110111111111111111110";
                        f_reg(161) <= "00000001110011010010000000100001";
                        f_reg(162) <= "00000011100110111001000000100001";
                        f_reg(163) <= "00000000100011000100000000100000";
                        f_reg(164) <= "00000010010110101011000000100000";
                        f_reg(165) <= "00000000000010110001101110000000";
                        f_reg(166) <= "00000000000110011000101110000000";
                        f_reg(167) <= "00000000001011010111000000100100";
                        f_reg(168) <= "00000001111110111110000000100100";
                        f_reg(169) <= "00000001010000100010000000100110";
                        f_reg(170) <= "00000011000100001001000000100110";
                        f_reg(171) <= "00000000000000000000000000000000";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00111100000010111000001101011100";
                        f_reg(174) <= "00111100000110011000001101011100";
                        f_reg(175) <= "00000000111010010000100000100100";
                        f_reg(176) <= "00000010101101110111100000100100";
                        f_reg(177) <= "00000001100011010101000000100010";
                        f_reg(178) <= "00000011010110111100000000100010";
                        f_reg(179) <= "10001100000001110000001111011000";
                        f_reg(180) <= "10001100000101010000001111011000";
                        f_reg(181) <= "00010100111101011111111111111110";
                        f_reg(182) <= "00000000111000110100100000000111";
                        f_reg(183) <= "00000010101100011011100000000111";
                        f_reg(184) <= "00000001001010000110000000100011";
                        f_reg(185) <= "00000010111101101101000000100011";
                        f_reg(186) <= "00010100101100110000000010101001";
                        f_reg(187) <= "10101100000001010000001110111000";
                        f_reg(188) <= "00000001010000010001100000100101";
                        f_reg(189) <= "00000011000011111000100000100101";
                        f_reg(190) <= "00010100011100010000000010100101";
                        f_reg(191) <= "10101100000000110000001110111100";
                        f_reg(192) <= "00000000000011000011100001000000";
                        f_reg(193) <= "00000000000110101010100001000000";
                        f_reg(194) <= "00110000110010011010011101011010";
                        f_reg(195) <= "00110010100101111010011101011010";
                        f_reg(196) <= "00000000100001110100000000000111";
                        f_reg(197) <= "00000010010101011011000000000111";
                        f_reg(198) <= "00000000000011100010110111000000";
                        f_reg(199) <= "00000000000111001001110111000000";
                        f_reg(200) <= "00000000010011010101000000101011";
                        f_reg(201) <= "00000010000110111100000000101011";
                        f_reg(202) <= "00000000101010000000100000000110";
                        f_reg(203) <= "00000010011101100111100000000110";
                        f_reg(204) <= "00100101011000110110000001101101";
                        f_reg(205) <= "00100111001100010110000001101101";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00010100011100010000000010001101";
                        f_reg(215) <= "10101100000000110000001111000000";
                        f_reg(216) <= "00010101010110000000000010001011";
                        f_reg(217) <= "10101100000010100000001111000100";
                        f_reg(218) <= "00010100010100000000000010001001";
                        f_reg(219) <= "10101100000000100000001111001000";
                        f_reg(220) <= "00010100001011110000000010000111";
                        f_reg(221) <= "10101100000000010000001111001100";
                        f_reg(222) <= "00010101001101110000000010000101";
                        f_reg(223) <= "10101100000010010000001111010000";
                        f_reg(224) <= "00100011110111011111111100000110";
                        f_reg(225) <= "00010011101000000000000000010111";
                        f_reg(226) <= "00100011110111011111111000001100";
                        f_reg(227) <= "00010011101000000000000000010101";
                        f_reg(228) <= "00100011110111011111110100010010";
                        f_reg(229) <= "00010011101000000000000000010011";
                        f_reg(230) <= "00100011110111101111111111111111";
                        f_reg(231) <= "00100011111111111111111111111111";
                        f_reg(232) <= "00010111110111110000000001111011";
                        f_reg(233) <= "00011111111000001111111101100101";
                        f_reg(234) <= "00010000000000000000000100000110";
                        f_reg(235) <= "00000000000000000000000000000000";
                        f_reg(236) <= "00000000000000000000000000000000";
                        f_reg(237) <= "00000000000000000000000000000000";
                        f_reg(238) <= "00000000000000000000000000000000";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000000000000000000000000000000";
                        f_reg(242) <= "00000000000000000000000000000000";
                        f_reg(243) <= "00000000000000000000000000000000";
                        f_reg(244) <= "00000000000000000000000000000000";
                        f_reg(245) <= "00000000000000000000000000000000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "10001100000111010000011100110000";
                        f_reg(249) <= "00011111101000000000000000000011";
                        f_reg(250) <= "00100000000111010000000000111100";
                        f_reg(251) <= "00010000000000000000000000000010";
                        f_reg(252) <= "00100000000111010000000000000000";
                        f_reg(253) <= "00010100001011110000000001100110";
                        f_reg(254) <= "10101111101000010000011010111000";
                        f_reg(255) <= "10001100000111010000011100110000";
                        f_reg(256) <= "00011111101000000000000000000011";
                        f_reg(257) <= "00100000000111010000000000111100";
                        f_reg(258) <= "00010000000000000000000000000010";
                        f_reg(259) <= "00100000000111010000000000000000";
                        f_reg(260) <= "00010100010100000000000001011111";
                        f_reg(261) <= "10101111101000100000011010111100";
                        f_reg(262) <= "10001100000111010000011100110000";
                        f_reg(263) <= "00011111101000000000000000000011";
                        f_reg(264) <= "00100000000111010000000000111100";
                        f_reg(265) <= "00010000000000000000000000000010";
                        f_reg(266) <= "00100000000111010000000000000000";
                        f_reg(267) <= "00010100011100010000000001011000";
                        f_reg(268) <= "10101111101000110000011011000000";
                        f_reg(269) <= "10001100000111010000011100110000";
                        f_reg(270) <= "00011111101000000000000000000011";
                        f_reg(271) <= "00100000000111010000000000111100";
                        f_reg(272) <= "00010000000000000000000000000010";
                        f_reg(273) <= "00100000000111010000000000000000";
                        f_reg(274) <= "00010100100100100000000001010001";
                        f_reg(275) <= "10101111101001000000011011000100";
                        f_reg(276) <= "10001100000111010000011100110000";
                        f_reg(277) <= "00011111101000000000000000000011";
                        f_reg(278) <= "00100000000111010000000000111100";
                        f_reg(279) <= "00010000000000000000000000000010";
                        f_reg(280) <= "00100000000111010000000000000000";
                        f_reg(281) <= "00010100101100110000000001001010";
                        f_reg(282) <= "10101111101001010000011011001000";
                        f_reg(283) <= "10001100000111010000011100110000";
                        f_reg(284) <= "00011111101000000000000000000011";
                        f_reg(285) <= "00100000000111010000000000111100";
                        f_reg(286) <= "00010000000000000000000000000010";
                        f_reg(287) <= "00100000000111010000000000000000";
                        f_reg(288) <= "00010100110101000000000001000011";
                        f_reg(289) <= "10101111101001100000011011001100";
                        f_reg(290) <= "10001100000111010000011100110000";
                        f_reg(291) <= "00011111101000000000000000000011";
                        f_reg(292) <= "00100000000111010000000000111100";
                        f_reg(293) <= "00010000000000000000000000000010";
                        f_reg(294) <= "00100000000111010000000000000000";
                        f_reg(295) <= "00010100111101010000000000111100";
                        f_reg(296) <= "10101111101001110000011011010000";
                        f_reg(297) <= "10001100000111010000011100110000";
                        f_reg(298) <= "00011111101000000000000000000011";
                        f_reg(299) <= "00100000000111010000000000111100";
                        f_reg(300) <= "00010000000000000000000000000010";
                        f_reg(301) <= "00100000000111010000000000000000";
                        f_reg(302) <= "00010101000101100000000000110101";
                        f_reg(303) <= "10101111101010000000011011010100";
                        f_reg(304) <= "10001100000111010000011100110000";
                        f_reg(305) <= "00011111101000000000000000000011";
                        f_reg(306) <= "00100000000111010000000000111100";
                        f_reg(307) <= "00010000000000000000000000000010";
                        f_reg(308) <= "00100000000111010000000000000000";
                        f_reg(309) <= "00010101001101110000000000101110";
                        f_reg(310) <= "10101111101010010000011011011000";
                        f_reg(311) <= "10001100000111010000011100110000";
                        f_reg(312) <= "00011111101000000000000000000011";
                        f_reg(313) <= "00100000000111010000000000111100";
                        f_reg(314) <= "00010000000000000000000000000010";
                        f_reg(315) <= "00100000000111010000000000000000";
                        f_reg(316) <= "00010101010110000000000000100111";
                        f_reg(317) <= "10101111101010100000011011011100";
                        f_reg(318) <= "10001100000111010000011100110000";
                        f_reg(319) <= "00011111101000000000000000000011";
                        f_reg(320) <= "00100000000111010000000000111100";
                        f_reg(321) <= "00010000000000000000000000000010";
                        f_reg(322) <= "00100000000111010000000000000000";
                        f_reg(323) <= "00010101011110010000000000100000";
                        f_reg(324) <= "10101111101010110000011011100000";
                        f_reg(325) <= "10001100000111010000011100110000";
                        f_reg(326) <= "00011111101000000000000000000011";
                        f_reg(327) <= "00100000000111010000000000111100";
                        f_reg(328) <= "00010000000000000000000000000010";
                        f_reg(329) <= "00100000000111010000000000000000";
                        f_reg(330) <= "00010101100110100000000000011001";
                        f_reg(331) <= "10101111101011000000011011100100";
                        f_reg(332) <= "10001100000111010000011100110000";
                        f_reg(333) <= "00011111101000000000000000000011";
                        f_reg(334) <= "00100000000111010000000000111100";
                        f_reg(335) <= "00010000000000000000000000000010";
                        f_reg(336) <= "00100000000111010000000000000000";
                        f_reg(337) <= "00010101101110110000000000010010";
                        f_reg(338) <= "10101111101011010000011011101000";
                        f_reg(339) <= "10001100000111010000011100110000";
                        f_reg(340) <= "00011111101000000000000000000011";
                        f_reg(341) <= "00100000000111010000000000111100";
                        f_reg(342) <= "00010000000000000000000000000010";
                        f_reg(343) <= "00100000000111010000000000000000";
                        f_reg(344) <= "00010101110111000000000000001011";
                        f_reg(345) <= "10101111101011100000011011101100";
                        f_reg(346) <= "10001100000111010000011100110000";
                        f_reg(347) <= "00011111101000000000000000000011";
                        f_reg(348) <= "00100000000111010000000000111100";
                        f_reg(349) <= "00010000000000000000000000000010";
                        f_reg(350) <= "00100000000111010000000000000000";
                        f_reg(351) <= "00010111110111110000000000000100";
                        f_reg(352) <= "10101111101111100000011011110000";
                        f_reg(353) <= "10101100000111010000011100110000";
                        f_reg(354) <= "00010000000000001111111110000100";
                        f_reg(355) <= "10001100000111010000011100110000";
                        f_reg(356) <= "10001111101000010000011010111000";
                        f_reg(357) <= "10001100000111010000011100110000";
                        f_reg(358) <= "10001111101011110000011010111000";
                        f_reg(359) <= "00010100001011111111111111111100";
                        f_reg(360) <= "10001100000111010000011100110000";
                        f_reg(361) <= "10001111101000100000011010111100";
                        f_reg(362) <= "10001100000111010000011100110000";
                        f_reg(363) <= "10001111101100000000011010111100";
                        f_reg(364) <= "00010100010100001111111111111100";
                        f_reg(365) <= "10001100000111010000011100110000";
                        f_reg(366) <= "10001111101000110000011011000000";
                        f_reg(367) <= "10001100000111010000011100110000";
                        f_reg(368) <= "10001111101100010000011011000000";
                        f_reg(369) <= "00010100011100011111111111111100";
                        f_reg(370) <= "10001100000111010000011100110000";
                        f_reg(371) <= "10001111101001000000011011000100";
                        f_reg(372) <= "10001100000111010000011100110000";
                        f_reg(373) <= "10001111101100100000011011000100";
                        f_reg(374) <= "00010100100100101111111111111100";
                        f_reg(375) <= "10001100000111010000011100110000";
                        f_reg(376) <= "10001111101001010000011011001000";
                        f_reg(377) <= "10001100000111010000011100110000";
                        f_reg(378) <= "10001111101100110000011011001000";
                        f_reg(379) <= "00010100101100111111111111111100";
                        f_reg(380) <= "10001100000111010000011100110000";
                        f_reg(381) <= "10001111101001100000011011001100";
                        f_reg(382) <= "10001100000111010000011100110000";
                        f_reg(383) <= "10001111101101000000011011001100";
                        f_reg(384) <= "00010100110101001111111111111100";
                        f_reg(385) <= "10001100000111010000011100110000";
                        f_reg(386) <= "10001111101001110000011011010000";
                        f_reg(387) <= "10001100000111010000011100110000";
                        f_reg(388) <= "10001111101101010000011011010000";
                        f_reg(389) <= "00010100111101011111111111111100";
                        f_reg(390) <= "10001100000111010000011100110000";
                        f_reg(391) <= "10001111101010000000011011010100";
                        f_reg(392) <= "10001100000111010000011100110000";
                        f_reg(393) <= "10001111101101100000011011010100";
                        f_reg(394) <= "00010101000101101111111111111100";
                        f_reg(395) <= "10001100000111010000011100110000";
                        f_reg(396) <= "10001111101010010000011011011000";
                        f_reg(397) <= "10001100000111010000011100110000";
                        f_reg(398) <= "10001111101101110000011011011000";
                        f_reg(399) <= "00010101001101111111111111111100";
                        f_reg(400) <= "10001100000111010000011100110000";
                        f_reg(401) <= "10001111101010100000011011011100";
                        f_reg(402) <= "10001100000111010000011100110000";
                        f_reg(403) <= "10001111101110000000011011011100";
                        f_reg(404) <= "00010101010110001111111111111100";
                        f_reg(405) <= "10001100000111010000011100110000";
                        f_reg(406) <= "10001111101010110000011011100000";
                        f_reg(407) <= "10001100000111010000011100110000";
                        f_reg(408) <= "10001111101110010000011011100000";
                        f_reg(409) <= "00010101011110011111111111111100";
                        f_reg(410) <= "10001100000111010000011100110000";
                        f_reg(411) <= "10001111101011000000011011100100";
                        f_reg(412) <= "10001100000111010000011100110000";
                        f_reg(413) <= "10001111101110100000011011100100";
                        f_reg(414) <= "00010101100110101111111111111100";
                        f_reg(415) <= "10001100000111010000011100110000";
                        f_reg(416) <= "10001111101011010000011011101000";
                        f_reg(417) <= "10001100000111010000011100110000";
                        f_reg(418) <= "10001111101110110000011011101000";
                        f_reg(419) <= "00010101101110111111111111111100";
                        f_reg(420) <= "10001100000111010000011100110000";
                        f_reg(421) <= "10001111101011100000011011101100";
                        f_reg(422) <= "10001100000111010000011100110000";
                        f_reg(423) <= "10001111101111000000011011101100";
                        f_reg(424) <= "00010101110111001111111111111100";
                        f_reg(425) <= "10001100000111010000011100110000";
                        f_reg(426) <= "10001111101111100000011011110000";
                        f_reg(427) <= "10001100000111010000011100110000";
                        f_reg(428) <= "10001111101111110000011011110000";
                        f_reg(429) <= "00010111110111111111111111111100";
                        f_reg(430) <= "00010000000000001111111100111000";
                        f_reg(431) <= "00000000000000000000000000000000";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000001111100111";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010011010011001001";
                        f_reg(4) <= "00111100000000101001011011000110";
                        f_reg(5) <= "00000000000000010001100000000110";
                        f_reg(6) <= "00101000001001000101110010010011";
                        f_reg(7) <= "10101100000001000000001110101000";
                        f_reg(8) <= "00000000000000000010100000100100";
                        f_reg(9) <= "00000000001000000011000000000110";
                        f_reg(10) <= "00000000110000010011100000100101";
                        f_reg(11) <= "00000000000000000000000000000000";
                        f_reg(12) <= "00000000110000000100000000100010";
                        f_reg(13) <= "00000000000010000100110101000000";
                        f_reg(14) <= "00100100101010101101000010011100";
                        f_reg(15) <= "00000001010001010101100000100011";
                        f_reg(16) <= "00101001011011000011010101010101";
                        f_reg(17) <= "00000000011001000110100000100110";
                        f_reg(18) <= "00000001100001100111000000101010";
                        f_reg(19) <= "00101001110011111011100100100011";
                        f_reg(20) <= "00000000001010111000000000000111";
                        f_reg(21) <= "10101100000010000000001110101100";
                        f_reg(22) <= "00000001101001111000100000000100";
                        f_reg(23) <= "00000000000000000000000000000000";
                        f_reg(24) <= "00000000010000011001000000100101";
                        f_reg(25) <= "00000001011011001001100000100010";
                        f_reg(26) <= "10101100000000100000001110110000";
                        f_reg(27) <= "00000001100011011010000000100101";
                        f_reg(28) <= "00000000000100111010111101000010";
                        f_reg(29) <= "00000010010001111011000000100100";
                        f_reg(30) <= "00110001001101110111010101110011";
                        f_reg(31) <= "00000000000011101100011011000011";
                        f_reg(32) <= "00000000010101011100100000000110";
                        f_reg(33) <= "00000010100001011101000000100011";
                        f_reg(34) <= "00111001110110111101011111110100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000000010100101110000000101010";
                        f_reg(37) <= "10101100000110100000001110110100";
                        f_reg(38) <= "00000010101101101110100000100000";
                        f_reg(39) <= "00000010001010001111000000100110";
                        f_reg(40) <= "00000010000110010101000000100101";
                        f_reg(41) <= "00000011100110000001100000100001";
                        f_reg(42) <= "00000000011010100010000000100000";
                        f_reg(43) <= "00000000000101000011001110000000";
                        f_reg(44) <= "00000010110110000000100000100100";
                        f_reg(45) <= "00000001111111010101100000100110";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00111100000011011000001101011100";
                        f_reg(48) <= "00000010111110011001100000100100";
                        f_reg(49) <= "00000001010110000011100000100010";
                        f_reg(50) <= "00000001100001100100100000000111";
                        f_reg(51) <= "00000001001001000010100000100011";
                        f_reg(52) <= "10101100000110110000001110111000";
                        f_reg(53) <= "00000000111100110111000000100101";
                        f_reg(54) <= "10101100000011100000001110111100";
                        f_reg(55) <= "00000000000001010001000001000000";
                        f_reg(56) <= "00110011110100101010011101011010";
                        f_reg(57) <= "00000001011000101101000000000111";
                        f_reg(58) <= "00000000000000011010110111000000";
                        f_reg(59) <= "00000011101110001000100000101011";
                        f_reg(60) <= "00000010101110100100000000000110";
                        f_reg(61) <= "00100101101100000110000001101101";
                        f_reg(62) <= "00000000000000000000000000000000";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000000000000000000000000000000";
                        f_reg(66) <= "10101100000100000000001111000000";
                        f_reg(67) <= "10101100000100010000001111000100";
                        f_reg(68) <= "10101100000111010000001111001000";
                        f_reg(69) <= "10101100000010000000001111001100";
                        f_reg(70) <= "10101100000100100000001111010000";
                        f_reg(71) <= "00100011111111111111111111111111";
                        f_reg(72) <= "00011111111000001111111110111011";
                        f_reg(73) <= "00010000000000000000000110100111";
                        f_reg(74) <= "00111100000111100000001111100111";
                        f_reg(75) <= "00111100000111110000001111100111";
                        f_reg(76) <= "00000000000111101111010000000010";
                        f_reg(77) <= "00000000000111111111110000000010";
                        f_reg(78) <= "00111100000000010011010011001001";
                        f_reg(79) <= "00111100000011110011010011001001";
                        f_reg(80) <= "00111100000000101001011011000110";
                        f_reg(81) <= "00111100000100001001011011000110";
                        f_reg(82) <= "00000000000000010001100000000110";
                        f_reg(83) <= "00000000000011111000100000000110";
                        f_reg(84) <= "00101000001001000101110010010011";
                        f_reg(85) <= "00101001111100100101110010010011";
                        f_reg(86) <= "00010100100100100000000100001101";
                        f_reg(87) <= "10101100000001000000001110101000";
                        f_reg(88) <= "00000000000000000010100000100100";
                        f_reg(89) <= "00000000000000001001100000100100";
                        f_reg(90) <= "00000000001000000011000000000110";
                        f_reg(91) <= "00000001111000001010000000000110";
                        f_reg(92) <= "00000000110000010011100000100101";
                        f_reg(93) <= "00000010100011111010100000100101";
                        f_reg(94) <= "00000000000000000000000000000000";
                        f_reg(95) <= "00000000000000000000000000000000";
                        f_reg(96) <= "00000000110000000100000000100010";
                        f_reg(97) <= "00000010100000001011000000100010";
                        f_reg(98) <= "00000000000010000100110101000000";
                        f_reg(99) <= "00000000000101101011110101000000";
                        f_reg(100) <= "00100100101010101101000010011100";
                        f_reg(101) <= "00100110011110001101000010011100";
                        f_reg(102) <= "00000001010001010101100000100011";
                        f_reg(103) <= "00000011000100111100100000100011";
                        f_reg(104) <= "00101001011011000011010101010101";
                        f_reg(105) <= "00101011001110100011010101010101";
                        f_reg(106) <= "00000000011001000110100000100110";
                        f_reg(107) <= "00000010001100101101100000100110";
                        f_reg(108) <= "00000001100001100111000000101010";
                        f_reg(109) <= "00000011010101001110000000101010";
                        f_reg(110) <= "00101001110010101011100100100011";
                        f_reg(111) <= "00101011100110001011100100100011";
                        f_reg(112) <= "00000000001010110001100000000111";
                        f_reg(113) <= "00000001111110011000100000000111";
                        f_reg(114) <= "00010101000101100000000011110001";
                        f_reg(115) <= "10101100000010000000001110101100";
                        f_reg(116) <= "00000001101001110010000000000100";
                        f_reg(117) <= "00000011011101011001000000000100";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000000000000000000000000000";
                        f_reg(120) <= "00000000010000010011000000100101";
                        f_reg(121) <= "00000010000011111010000000100101";
                        f_reg(122) <= "00000001011011000000100000100010";
                        f_reg(123) <= "00000011001110100111100000100010";
                        f_reg(124) <= "00010100010100000000000011100111";
                        f_reg(125) <= "10101100000000100000001110110000";
                        f_reg(126) <= "00000001100011010101100000100101";
                        f_reg(127) <= "00000011010110111100100000100101";
                        f_reg(128) <= "00000000000000010110111101000010";
                        f_reg(129) <= "00000000000011111101111101000010";
                        f_reg(130) <= "00000000110001110000100000100100";
                        f_reg(131) <= "00000010100101010111100000100100";
                        f_reg(132) <= "00110001001001110111010101110011";
                        f_reg(133) <= "00110010111101010111010101110011";
                        f_reg(134) <= "00000000000011100100111011000011";
                        f_reg(135) <= "00000000000111001011111011000011";
                        f_reg(136) <= "00010101001101110000000011011011";
                        f_reg(137) <= "10101100000010010000001111010100";
                        f_reg(138) <= "00000000010011010100100000000110";
                        f_reg(139) <= "00000010000110111011100000000110";
                        f_reg(140) <= "00010101100110100000000011010111";
                        f_reg(141) <= "10101100000011000000001111011000";
                        f_reg(142) <= "00000001011001010110000000100011";
                        f_reg(143) <= "00000011001100111101000000100011";
                        f_reg(144) <= "00111001110001011101011111110100";
                        f_reg(145) <= "00111011100100111101011111110100";
                        f_reg(146) <= "00000000000000000000000000000000";
                        f_reg(147) <= "00000000000000000000000000000000";
                        f_reg(148) <= "00000000010001100111000000101010";
                        f_reg(149) <= "00000010000101001110000000101010";
                        f_reg(150) <= "00010101100110100000000011001101";
                        f_reg(151) <= "10101100000011000000001110110100";
                        f_reg(152) <= "00000001101000010001000000100000";
                        f_reg(153) <= "00000011011011111000000000100000";
                        f_reg(154) <= "00000000100010000011000000100110";
                        f_reg(155) <= "00000010010101101010000000100110";
                        f_reg(156) <= "00000000011010010110000000100101";
                        f_reg(157) <= "00000010001101111101000000100101";
                        f_reg(158) <= "10001100000011010000001111010100";
                        f_reg(159) <= "10001100000110110000001111010100";
                        f_reg(160) <= "00010101101110111111111111111110";
                        f_reg(161) <= "00000001110011010010000000100001";
                        f_reg(162) <= "00000011100110111001000000100001";
                        f_reg(163) <= "00000000100011000100000000100000";
                        f_reg(164) <= "00000010010110101011000000100000";
                        f_reg(165) <= "00000000000010110001101110000000";
                        f_reg(166) <= "00000000000110011000101110000000";
                        f_reg(167) <= "00000000001011010111000000100100";
                        f_reg(168) <= "00000001111110111110000000100100";
                        f_reg(169) <= "00000001010000100010000000100110";
                        f_reg(170) <= "00000011000100001001000000100110";
                        f_reg(171) <= "00000000000000000000000000000000";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00111100000010111000001101011100";
                        f_reg(174) <= "00111100000110011000001101011100";
                        f_reg(175) <= "00000000111010010000100000100100";
                        f_reg(176) <= "00000010101101110111100000100100";
                        f_reg(177) <= "00000001100011010101000000100010";
                        f_reg(178) <= "00000011010110111100000000100010";
                        f_reg(179) <= "10001100000001110000001111011000";
                        f_reg(180) <= "10001100000101010000001111011000";
                        f_reg(181) <= "00010100111101011111111111111110";
                        f_reg(182) <= "00000000111000110100100000000111";
                        f_reg(183) <= "00000010101100011011100000000111";
                        f_reg(184) <= "00000001001010000110000000100011";
                        f_reg(185) <= "00000010111101101101000000100011";
                        f_reg(186) <= "00010100101100110000000010101001";
                        f_reg(187) <= "10101100000001010000001110111000";
                        f_reg(188) <= "00000001010000010001100000100101";
                        f_reg(189) <= "00000011000011111000100000100101";
                        f_reg(190) <= "00010100011100010000000010100101";
                        f_reg(191) <= "10101100000000110000001110111100";
                        f_reg(192) <= "00000000000011000011100001000000";
                        f_reg(193) <= "00000000000110101010100001000000";
                        f_reg(194) <= "00110000110010011010011101011010";
                        f_reg(195) <= "00110010100101111010011101011010";
                        f_reg(196) <= "00000000100001110100000000000111";
                        f_reg(197) <= "00000010010101011011000000000111";
                        f_reg(198) <= "00000000000011100010110111000000";
                        f_reg(199) <= "00000000000111001001110111000000";
                        f_reg(200) <= "00000000010011010101000000101011";
                        f_reg(201) <= "00000010000110111100000000101011";
                        f_reg(202) <= "00000000101010000000100000000110";
                        f_reg(203) <= "00000010011101100111100000000110";
                        f_reg(204) <= "00100101011000110110000001101101";
                        f_reg(205) <= "00100111001100010110000001101101";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00010100011100010000000010001101";
                        f_reg(215) <= "10101100000000110000001111000000";
                        f_reg(216) <= "00010101010110000000000010001011";
                        f_reg(217) <= "10101100000010100000001111000100";
                        f_reg(218) <= "00010100010100000000000010001001";
                        f_reg(219) <= "10101100000000100000001111001000";
                        f_reg(220) <= "00010100001011110000000010000111";
                        f_reg(221) <= "10101100000000010000001111001100";
                        f_reg(222) <= "00010101001101110000000010000101";
                        f_reg(223) <= "10101100000010010000001111010000";
                        f_reg(224) <= "00100011110111011111111100000110";
                        f_reg(225) <= "00010011101000000000000000010111";
                        f_reg(226) <= "00100011110111011111111000001100";
                        f_reg(227) <= "00010011101000000000000000010101";
                        f_reg(228) <= "00100011110111011111110100010010";
                        f_reg(229) <= "00010011101000000000000000010011";
                        f_reg(230) <= "00100011110111101111111111111111";
                        f_reg(231) <= "00100011111111111111111111111111";
                        f_reg(232) <= "00010111110111110000000001111011";
                        f_reg(233) <= "00011111111000001111111101100101";
                        f_reg(234) <= "00010000000000000000000100000110";
                        f_reg(235) <= "00000000000000000000000000000000";
                        f_reg(236) <= "00000000000000000000000000000000";
                        f_reg(237) <= "00000000000000000000000000000000";
                        f_reg(238) <= "00000000000000000000000000000000";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000000000000000000000000000000";
                        f_reg(242) <= "00000000000000000000000000000000";
                        f_reg(243) <= "00000000000000000000000000000000";
                        f_reg(244) <= "00000000000000000000000000000000";
                        f_reg(245) <= "00000000000000000000000000000000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "10001100000111010000011100110000";
                        f_reg(249) <= "00011111101000000000000000000011";
                        f_reg(250) <= "00100000000111010000000000111100";
                        f_reg(251) <= "00010000000000000000000000000010";
                        f_reg(252) <= "00100000000111010000000000000000";
                        f_reg(253) <= "00010100001011110000000001100110";
                        f_reg(254) <= "10101111101000010000011010111000";
                        f_reg(255) <= "10001100000111010000011100110000";
                        f_reg(256) <= "00011111101000000000000000000011";
                        f_reg(257) <= "00100000000111010000000000111100";
                        f_reg(258) <= "00010000000000000000000000000010";
                        f_reg(259) <= "00100000000111010000000000000000";
                        f_reg(260) <= "00010100010100000000000001011111";
                        f_reg(261) <= "10101111101000100000011010111100";
                        f_reg(262) <= "10001100000111010000011100110000";
                        f_reg(263) <= "00011111101000000000000000000011";
                        f_reg(264) <= "00100000000111010000000000111100";
                        f_reg(265) <= "00010000000000000000000000000010";
                        f_reg(266) <= "00100000000111010000000000000000";
                        f_reg(267) <= "00010100011100010000000001011000";
                        f_reg(268) <= "10101111101000110000011011000000";
                        f_reg(269) <= "10001100000111010000011100110000";
                        f_reg(270) <= "00011111101000000000000000000011";
                        f_reg(271) <= "00100000000111010000000000111100";
                        f_reg(272) <= "00010000000000000000000000000010";
                        f_reg(273) <= "00100000000111010000000000000000";
                        f_reg(274) <= "00010100100100100000000001010001";
                        f_reg(275) <= "10101111101001000000011011000100";
                        f_reg(276) <= "10001100000111010000011100110000";
                        f_reg(277) <= "00011111101000000000000000000011";
                        f_reg(278) <= "00100000000111010000000000111100";
                        f_reg(279) <= "00010000000000000000000000000010";
                        f_reg(280) <= "00100000000111010000000000000000";
                        f_reg(281) <= "00010100101100110000000001001010";
                        f_reg(282) <= "10101111101001010000011011001000";
                        f_reg(283) <= "10001100000111010000011100110000";
                        f_reg(284) <= "00011111101000000000000000000011";
                        f_reg(285) <= "00100000000111010000000000111100";
                        f_reg(286) <= "00010000000000000000000000000010";
                        f_reg(287) <= "00100000000111010000000000000000";
                        f_reg(288) <= "00010100110101000000000001000011";
                        f_reg(289) <= "10101111101001100000011011001100";
                        f_reg(290) <= "10001100000111010000011100110000";
                        f_reg(291) <= "00011111101000000000000000000011";
                        f_reg(292) <= "00100000000111010000000000111100";
                        f_reg(293) <= "00010000000000000000000000000010";
                        f_reg(294) <= "00100000000111010000000000000000";
                        f_reg(295) <= "00010100111101010000000000111100";
                        f_reg(296) <= "10101111101001110000011011010000";
                        f_reg(297) <= "10001100000111010000011100110000";
                        f_reg(298) <= "00011111101000000000000000000011";
                        f_reg(299) <= "00100000000111010000000000111100";
                        f_reg(300) <= "00010000000000000000000000000010";
                        f_reg(301) <= "00100000000111010000000000000000";
                        f_reg(302) <= "00010101000101100000000000110101";
                        f_reg(303) <= "10101111101010000000011011010100";
                        f_reg(304) <= "10001100000111010000011100110000";
                        f_reg(305) <= "00011111101000000000000000000011";
                        f_reg(306) <= "00100000000111010000000000111100";
                        f_reg(307) <= "00010000000000000000000000000010";
                        f_reg(308) <= "00100000000111010000000000000000";
                        f_reg(309) <= "00010101001101110000000000101110";
                        f_reg(310) <= "10101111101010010000011011011000";
                        f_reg(311) <= "10001100000111010000011100110000";
                        f_reg(312) <= "00011111101000000000000000000011";
                        f_reg(313) <= "00100000000111010000000000111100";
                        f_reg(314) <= "00010000000000000000000000000010";
                        f_reg(315) <= "00100000000111010000000000000000";
                        f_reg(316) <= "00010101010110000000000000100111";
                        f_reg(317) <= "10101111101010100000011011011100";
                        f_reg(318) <= "10001100000111010000011100110000";
                        f_reg(319) <= "00011111101000000000000000000011";
                        f_reg(320) <= "00100000000111010000000000111100";
                        f_reg(321) <= "00010000000000000000000000000010";
                        f_reg(322) <= "00100000000111010000000000000000";
                        f_reg(323) <= "00010101011110010000000000100000";
                        f_reg(324) <= "10101111101010110000011011100000";
                        f_reg(325) <= "10001100000111010000011100110000";
                        f_reg(326) <= "00011111101000000000000000000011";
                        f_reg(327) <= "00100000000111010000000000111100";
                        f_reg(328) <= "00010000000000000000000000000010";
                        f_reg(329) <= "00100000000111010000000000000000";
                        f_reg(330) <= "00010101100110100000000000011001";
                        f_reg(331) <= "10101111101011000000011011100100";
                        f_reg(332) <= "10001100000111010000011100110000";
                        f_reg(333) <= "00011111101000000000000000000011";
                        f_reg(334) <= "00100000000111010000000000111100";
                        f_reg(335) <= "00010000000000000000000000000010";
                        f_reg(336) <= "00100000000111010000000000000000";
                        f_reg(337) <= "00010101101110110000000000010010";
                        f_reg(338) <= "10101111101011010000011011101000";
                        f_reg(339) <= "10001100000111010000011100110000";
                        f_reg(340) <= "00011111101000000000000000000011";
                        f_reg(341) <= "00100000000111010000000000111100";
                        f_reg(342) <= "00010000000000000000000000000010";
                        f_reg(343) <= "00100000000111010000000000000000";
                        f_reg(344) <= "00010101110111000000000000001011";
                        f_reg(345) <= "10101111101011100000011011101100";
                        f_reg(346) <= "10001100000111010000011100110000";
                        f_reg(347) <= "00011111101000000000000000000011";
                        f_reg(348) <= "00100000000111010000000000111100";
                        f_reg(349) <= "00010000000000000000000000000010";
                        f_reg(350) <= "00100000000111010000000000000000";
                        f_reg(351) <= "00010111110111110000000000000100";
                        f_reg(352) <= "10101111101111100000011011110000";
                        f_reg(353) <= "10101100000111010000011100110000";
                        f_reg(354) <= "00010000000000001111111110000100";
                        f_reg(355) <= "10001100000111010000011100110000";
                        f_reg(356) <= "10001111101000010000011010111000";
                        f_reg(357) <= "10001100000111010000011100110000";
                        f_reg(358) <= "10001111101011110000011010111000";
                        f_reg(359) <= "00010100001011111111111111111100";
                        f_reg(360) <= "10001100000111010000011100110000";
                        f_reg(361) <= "10001111101000100000011010111100";
                        f_reg(362) <= "10001100000111010000011100110000";
                        f_reg(363) <= "10001111101100000000011010111100";
                        f_reg(364) <= "00010100010100001111111111111100";
                        f_reg(365) <= "10001100000111010000011100110000";
                        f_reg(366) <= "10001111101000110000011011000000";
                        f_reg(367) <= "10001100000111010000011100110000";
                        f_reg(368) <= "10001111101100010000011011000000";
                        f_reg(369) <= "00010100011100011111111111111100";
                        f_reg(370) <= "10001100000111010000011100110000";
                        f_reg(371) <= "10001111101001000000011011000100";
                        f_reg(372) <= "10001100000111010000011100110000";
                        f_reg(373) <= "10001111101100100000011011000100";
                        f_reg(374) <= "00010100100100101111111111111100";
                        f_reg(375) <= "10001100000111010000011100110000";
                        f_reg(376) <= "10001111101001010000011011001000";
                        f_reg(377) <= "10001100000111010000011100110000";
                        f_reg(378) <= "10001111101100110000011011001000";
                        f_reg(379) <= "00010100101100111111111111111100";
                        f_reg(380) <= "10001100000111010000011100110000";
                        f_reg(381) <= "10001111101001100000011011001100";
                        f_reg(382) <= "10001100000111010000011100110000";
                        f_reg(383) <= "10001111101101000000011011001100";
                        f_reg(384) <= "00010100110101001111111111111100";
                        f_reg(385) <= "10001100000111010000011100110000";
                        f_reg(386) <= "10001111101001110000011011010000";
                        f_reg(387) <= "10001100000111010000011100110000";
                        f_reg(388) <= "10001111101101010000011011010000";
                        f_reg(389) <= "00010100111101011111111111111100";
                        f_reg(390) <= "10001100000111010000011100110000";
                        f_reg(391) <= "10001111101010000000011011010100";
                        f_reg(392) <= "10001100000111010000011100110000";
                        f_reg(393) <= "10001111101101100000011011010100";
                        f_reg(394) <= "00010101000101101111111111111100";
                        f_reg(395) <= "10001100000111010000011100110000";
                        f_reg(396) <= "10001111101010010000011011011000";
                        f_reg(397) <= "10001100000111010000011100110000";
                        f_reg(398) <= "10001111101101110000011011011000";
                        f_reg(399) <= "00010101001101111111111111111100";
                        f_reg(400) <= "10001100000111010000011100110000";
                        f_reg(401) <= "10001111101010100000011011011100";
                        f_reg(402) <= "10001100000111010000011100110000";
                        f_reg(403) <= "10001111101110000000011011011100";
                        f_reg(404) <= "00010101010110001111111111111100";
                        f_reg(405) <= "10001100000111010000011100110000";
                        f_reg(406) <= "10001111101010110000011011100000";
                        f_reg(407) <= "10001100000111010000011100110000";
                        f_reg(408) <= "10001111101110010000011011100000";
                        f_reg(409) <= "00010101011110011111111111111100";
                        f_reg(410) <= "10001100000111010000011100110000";
                        f_reg(411) <= "10001111101011000000011011100100";
                        f_reg(412) <= "10001100000111010000011100110000";
                        f_reg(413) <= "10001111101110100000011011100100";
                        f_reg(414) <= "00010101100110101111111111111100";
                        f_reg(415) <= "10001100000111010000011100110000";
                        f_reg(416) <= "10001111101011010000011011101000";
                        f_reg(417) <= "10001100000111010000011100110000";
                        f_reg(418) <= "10001111101110110000011011101000";
                        f_reg(419) <= "00010101101110111111111111111100";
                        f_reg(420) <= "10001100000111010000011100110000";
                        f_reg(421) <= "10001111101011100000011011101100";
                        f_reg(422) <= "10001100000111010000011100110000";
                        f_reg(423) <= "10001111101111000000011011101100";
                        f_reg(424) <= "00010101110111001111111111111100";
                        f_reg(425) <= "10001100000111010000011100110000";
                        f_reg(426) <= "10001111101111100000011011110000";
                        f_reg(427) <= "10001100000111010000011100110000";
                        f_reg(428) <= "10001111101111110000011011110000";
                        f_reg(429) <= "00010111110111111111111111111100";
                        f_reg(430) <= "00010000000000001111111100111000";
                        f_reg(431) <= "00000000000000000000000000000000";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000001111100111";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test73_Reg_COMBINED;
