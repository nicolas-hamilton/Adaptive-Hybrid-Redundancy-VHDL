--| Test20_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:09:23
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test20_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test20_Reg_COMBINED;

architecture a_Test20_Reg_COMBINED of Test20_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 540) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 540) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100", --  495 - 1980
      "00000000000000000000011111000000", --  496 - 1984
      "00000000000000000000011111000100", --  497 - 1988
      "00000000000000000000011111001000", --  498 - 1992
      "00000000000000000000011111001100", --  499 - 1996
      "00000000000000000000011111010000", --  500 - 2000
      "00000000000000000000011111010100", --  501 - 2004
      "00000000000000000000011111011000", --  502 - 2008
      "00000000000000000000011111011100", --  503 - 2012
      "00000000000000000000011111100000", --  504 - 2016
      "00000000000000000000011111100100", --  505 - 2020
      "00000000000000000000011111101000", --  506 - 2024
      "00000000000000000000011111101100", --  507 - 2028
      "00000000000000000000011111110000", --  508 - 2032
      "00000000000000000000011111110100", --  509 - 2036
      "00000000000000000000011111111000", --  510 - 2040
      "00000000000000000000011111111100", --  511 - 2044
      "00000000000000000000100000000000", --  512 - 2048
      "00000000000000000000100000000100", --  513 - 2052
      "00000000000000000000100000001000", --  514 - 2056
      "00000000000000000000100000001100", --  515 - 2060
      "00000000000000000000100000010000", --  516 - 2064
      "00000000000000000000100000010100", --  517 - 2068
      "00000000000000000000100000011000", --  518 - 2072
      "00000000000000000000100000011100", --  519 - 2076
      "00000000000000000000100000100000", --  520 - 2080
      "00000000000000000000100000100100", --  521 - 2084
      "00000000000000000000100000101000", --  522 - 2088
      "00000000000000000000100000101100", --  523 - 2092
      "00000000000000000000100000110000", --  524 - 2096
      "00000000000000000000100000110100", --  525 - 2100
      "00000000000000000000100000111000", --  526 - 2104
      "00000000000000000000100000111100", --  527 - 2108
      "00000000000000000000100001000000", --  528 - 2112
      "00000000000000000000100001000100", --  529 - 2116
      "00000000000000000000100001001000", --  530 - 2120
      "00000000000000000000100001001100", --  531 - 2124
      "00000000000000000000100001010000", --  532 - 2128
      "00000000000000000000100001010100", --  533 - 2132
      "00000000000000000000100001011000", --  534 - 2136
      "00000000000000000000100001011100", --  535 - 2140
      "00000000000000000000100001100000", --  536 - 2144
      "00000000000000000000100001100100", --  537 - 2148
      "00000000000000000000100001101000", --  538 - 2152
      "00000000000000000000100001101100");--  539 - 2156

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000010001001011010101", --    2 -    8
      "00000000001000010001000000100010", --    3 -   12
      "00101000001000110010100010011111", --    4 -   16
      "00000000001000010010000000100000", --    5 -   20
      "00000000000000100010100001000011", --    6 -   24
      "00000000101000110011000000100011", --    7 -   28
      "00000000010000100011100000100101", --    8 -   32
      "00000000000000000100000111000011", --    9 -   36
      "10101100000010000000010001000000", --   10 -   40
      "10101100000000010000010001000100", --   11 -   44
      "00000000100001000100100000000110", --   12 -   48
      "00000000111001110101000000101011", --   13 -   52
      "00000000110010100101100000100111", --   14 -   56
      "10101100000010000000010001001000", --   15 -   60
      "00000001000000010110000000000100", --   16 -   64
      "00000000000000000000000000000000", --   17 -   68
      "00000001100010110110100000101011", --   18 -   72
      "00000000000010000111000110000010", --   19 -   76
      "10101100000000010000010001001100", --   20 -   80
      "00000001001001010010100000101011", --   21 -   84
      "00000000001001100111100000100011", --   22 -   88
      "00000000100000111000000000100100", --   23 -   92
      "00101001110100011000100100101101", --   24 -   96
      "00000000100001101001000000100111", --   25 -  100
      "00101101000100110100100000000010", --   26 -  104
      "00000001101000011010000000100100", --   27 -  108
      "10101100000011000000010001010000", --   28 -  112
      "00000000000000011010100000000110", --   29 -  116
      "00000010010011101011000000100001", --   30 -  120
      "00000000101011111011100000101010", --   31 -  124
      "00000001011010101100000000100001", --   32 -  128
      "10101100000010100000010001010100", --   33 -  132
      "00000000000000000000000000000000", --   34 -  136
      "00000010011100101100100000100101", --   35 -  140
      "00000000000010011101010000000011", --   36 -  144
      "10101100000110010000010001011000", --   37 -  148
      "00000000110001000011000000100010", --   38 -  152
      "00100110111110111101010011110111", --   39 -  156
      "00000000101011010010100000100111", --   40 -  160
      "00000000000110011110010000000011", --   41 -  164
      "00101101011111010001011001001101", --   42 -  168
      "00000011011100001111000000101011", --   43 -  172
      "00000011000100100001000000100000", --   44 -  176
      "00000010100000000011100000100100", --   45 -  180
      "10101100000001110000010001011100", --   46 -  184
      "00110010101000111000000001111000", --   47 -  188
      "00000000010111100110000000100011", --   48 -  192
      "00000011010111000000100000100010", --   49 -  196
      "00000000110111100111000000101011", --   50 -  200
      "00000000010010000111100000100101", --   51 -  204
      "00100111001010101000000100111100", --   52 -  208
      "00111000101010011100000101001101", --   53 -  212
      "10101100000100010000010001100000", --   54 -  216
      "00101101110001000110110111011111", --   55 -  220
      "10101100000011110000010001100100", --   56 -  224
      "10101100000010100000010001101000", --   57 -  228
      "00000011110010011011100000000100", --   58 -  232
      "00000000011111010110100000101010", --   59 -  236
      "00000000001001000101100000100110", --   60 -  240
      "00000000110011101101100000100111", --   61 -  244
      "00000000000000000000000000000000", --   62 -  248
      "10101100000110110000010001101100", --   63 -  252
      "10101100000011010000010001110000", --   64 -  256
      "00000010111000001000000000100100", --   65 -  260
      "00000010011011001100000000100010", --   66 -  264
      "00000010110010111001000000100000", --   67 -  268
      "00000000000000000000000000000000", --   68 -  272
      "00110110000101000111000001000101", --   69 -  276
      "00000000000000000000000000000000", --   70 -  280
      "00000010100110000011100000101011", --   71 -  284
      "10101100000001110000010001110100", --   72 -  288
      "00000000000100101001001111000000", --   73 -  292
      "00000000000000000000000000000000", --   74 -  296
      "10101100000100100000010001111000", --   75 -  300
      "00100011111111111111111111111111", --   76 -  304
      "00011111111000001111111110110101", --   77 -  308
      "00010000000000000000000111001101", --   78 -  312
      "00111100000111100000001111100111", --   79 -  316
      "00111100000111110000001111100111", --   80 -  320
      "00000000000111101111010000000010", --   81 -  324
      "00000000000111111111110000000010", --   82 -  328
      "00111100000000010001001011010101", --   83 -  332
      "00111100000011110001001011010101", --   84 -  336
      "00000000001000010001000000100010", --   85 -  340
      "00000001111011111000000000100010", --   86 -  344
      "00101000001000110010100010011111", --   87 -  348
      "00101001111100010010100010011111", --   88 -  352
      "00000000001000010010000000100000", --   89 -  356
      "00000001111011111001000000100000", --   90 -  360
      "00000000000000100010100001000011", --   91 -  364
      "00000000000100001001100001000011", --   92 -  368
      "00000000101000110011000000100011", --   93 -  372
      "00000010011100011010000000100011", --   94 -  376
      "00000000010000100011100000100101", --   95 -  380
      "00000010000100001010100000100101", --   96 -  384
      "00000000000000000100000111000011", --   97 -  388
      "00000000000000001011000111000011", --   98 -  392
      "00010101000101100000000100101011", --   99 -  396
      "10101100000010000000010001000000", --  100 -  400
      "00010100001011110000000100101001", --  101 -  404
      "10101100000000010000010001000100", --  102 -  408
      "00000000100001000100100000000110", --  103 -  412
      "00000010010100101011100000000110", --  104 -  416
      "00000000111001110101000000101011", --  105 -  420
      "00000010101101011100000000101011", --  106 -  424
      "00000000110010100101100000100111", --  107 -  428
      "00000010100110001100100000100111", --  108 -  432
      "00010101000101100000000100100001", --  109 -  436
      "10101100000010000000010001001000", --  110 -  440
      "00000001000000010110000000000100", --  111 -  444
      "00000010110011111101000000000100", --  112 -  448
      "00000000000000000000000000000000", --  113 -  452
      "00000000000000000000000000000000", --  114 -  456
      "00000001100010110110100000101011", --  115 -  460
      "00000011010110011101100000101011", --  116 -  464
      "00000000000010000111000110000010", --  117 -  468
      "00000000000101101110000110000010", --  118 -  472
      "00010100001011110000000100010111", --  119 -  476
      "10101100000000010000010001001100", --  120 -  480
      "00000001001001010010100000101011", --  121 -  484
      "00000010111100111001100000101011", --  122 -  488
      "00000000001001100001000000100011", --  123 -  492
      "00000001111101001000000000100011", --  124 -  496
      "00000000100000110011100000100100", --  125 -  500
      "00000010010100011010100000100100", --  126 -  504
      "00101001110000111000100100101101", --  127 -  508
      "00101011100100011000100100101101", --  128 -  512
      "00010100011100010000000100001101", --  129 -  516
      "10101100000000110000010001111100", --  130 -  520
      "00000000100001100001100000100111", --  131 -  524
      "00000010010101001000100000100111", --  132 -  528
      "00010100011100010000000100001001", --  133 -  532
      "10101100000000110000010010000000", --  134 -  536
      "00101101000000110100100000000010", --  135 -  540
      "00101110110100010100100000000010", --  136 -  544
      "00010100011100010000000100000101", --  137 -  548
      "10101100000000110000010010000100", --  138 -  552
      "00000001101000010001100000100100", --  139 -  556
      "00000011011011111000100000100100", --  140 -  560
      "00010101100110100000000100000001", --  141 -  564
      "10101100000011000000010001010000", --  142 -  568
      "00000000000000010110000000000110", --  143 -  572
      "00000000000011111101000000000110", --  144 -  576
      "10001100000000010000010010000000", --  145 -  580
      "10001100000011110000010010000000", --  146 -  584
      "00010100001011111111111111111110", --  147 -  588
      "00010101000101100000000011111010", --  148 -  592
      "10101100000010000000010010000000", --  149 -  596
      "00000000001011100100000000100001", --  150 -  600
      "00000001111111001011000000100001", --  151 -  604
      "00000000101000100111000000101010", --  152 -  608
      "00000010011100001110000000101010", --  153 -  612
      "00000001011010100001000000100001", --  154 -  616
      "00000011001110001000000000100001", --  155 -  620
      "00010101010110000000000011110010", --  156 -  624
      "10101100000010100000010001010100", --  157 -  628
      "00000000000000000000000000000000", --  158 -  632
      "00000000000000000000000000000000", --  159 -  636
      "10001100000010100000010010000100", --  160 -  640
      "10001100000110000000010010000100", --  161 -  644
      "00010101010110001111111111111110", --  162 -  648
      "00010101000101100000000011101011", --  163 -  652
      "10101100000010000000010010000100", --  164 -  656
      "00000001010000010100000000100101", --  165 -  660
      "00000011000011111011000000100101", --  166 -  664
      "00010101010110000000000011100111", --  167 -  668
      "10101100000010100000010010001000", --  168 -  672
      "00000000000010010101010000000011", --  169 -  676
      "00000000000101111100010000000011", --  170 -  680
      "00010101000101100000000011100011", --  171 -  684
      "10101100000010000000010001011000", --  172 -  688
      "00000000110001000011000000100010", --  173 -  692
      "00000010100100101010000000100010", --  174 -  696
      "00100101110010011101010011110111", --  175 -  700
      "00100111100101111101010011110111", --  176 -  704
      "00000000101011010010100000100111", --  177 -  708
      "00000010011110111001100000100111", --  178 -  712
      "00000000000010000010010000000011", --  179 -  716
      "00000000000101101001010000000011", --  180 -  720
      "00101101011011100001011001001101", --  181 -  724
      "00101111001111000001011001001101", --  182 -  728
      "00000001001001110110100000101011", --  183 -  732
      "00000010111101011101100000101011", --  184 -  736
      "00000000010000010101100000100000", --  185 -  740
      "00000010000011111100100000100000", --  186 -  744
      "00000000011000000100100000100100", --  187 -  748
      "00000010001000001011100000100100", --  188 -  752
      "00010101001101110000000011010001", --  189 -  756
      "10101100000010010000010001011100", --  190 -  760
      "00110001100001111000000001111000", --  191 -  764
      "00110011010101011000000001111000", --  192 -  768
      "00000001011011010001000000100011", --  193 -  772
      "00000011001110111000000000100011", --  194 -  776
      "00000001010001000000100000100010", --  195 -  780
      "00000011000100100111100000100010", --  196 -  784
      "00000000110011010001100000101011", --  197 -  788
      "00000010100110111000100000101011", --  198 -  792
      "10001100000010010000010010000000", --  199 -  796
      "10001100000101110000010010000000", --  200 -  800
      "00010101001101111111111111111110", --  201 -  804
      "00000001011010010110000000100101", --  202 -  808
      "00000011001101111101000000100101", --  203 -  812
      "00100101000010101000000100111100", --  204 -  816
      "00100110110110001000000100111100", --  205 -  820
      "00111000101001001100000101001101", --  206 -  824
      "00111010011100101100000101001101", --  207 -  828
      "10001100000010110000010001111100", --  208 -  832
      "10001100000110010000010001111100", --  209 -  836
      "00010101011110011111111111111110", --  210 -  840
      "00010101011110010000000010111011", --  211 -  844
      "10101100000010110000010001100000", --  212 -  848
      "00101100011010010110110111011111", --  213 -  852
      "00101110001101110110110111011111", --  214 -  856
      "00010101100110100000000010110111", --  215 -  860
      "10101100000011000000010001100100", --  216 -  864
      "00010101010110000000000010110101", --  217 -  868
      "10101100000010100000010001101000", --  218 -  872
      "00000001101001000100000000000100", --  219 -  876
      "00000011011100101011000000000100", --  220 -  880
      "00000000111011100010100000101010", --  221 -  884
      "00000010101111001001100000101010", --  222 -  888
      "00000000001010010101100000100110", --  223 -  892
      "00000001111101111100100000100110", --  224 -  896
      "00000000110000110110000000100111", --  225 -  900
      "00000010100100011101000000100111", --  226 -  904
      "00000000000000000000000000000000", --  227 -  908
      "00000000000000000000000000000000", --  228 -  912
      "00010101100110100000000010101001", --  229 -  916
      "10101100000011000000010001101100", --  230 -  920
      "00010100101100110000000010100111", --  231 -  924
      "10101100000001010000010001110000", --  232 -  928
      "00000001000000000101000000100100", --  233 -  932
      "00000010110000001100000000100100", --  234 -  936
      "10001100000001000000010010001000", --  235 -  940
      "10001100000100100000010010001000", --  236 -  944
      "00010100100100101111111111111110", --  237 -  948
      "00000000100000100110100000100010", --  238 -  952
      "00000010010100001101100000100010", --  239 -  956
      "10001100000001110000010010000100", --  240 -  960
      "10001100000101010000010010000100", --  241 -  964
      "00010100111101011111111111111110", --  242 -  968
      "00000000111010110111000000100000", --  243 -  972
      "00000010101110011110000000100000", --  244 -  976
      "00000000000000000000000000000000", --  245 -  980
      "00000000000000000000000000000000", --  246 -  984
      "00110101010000010111000001000101", --  247 -  988
      "00110111000011110111000001000101", --  248 -  992
      "00000000000000000000000000000000", --  249 -  996
      "00000000000000000000000000000000", --  250 - 1000
      "00000000001011010100100000101011", --  251 - 1004
      "00000001111110111011100000101011", --  252 - 1008
      "00010101001101110000000010010001", --  253 - 1012
      "10101100000010010000010001110100", --  254 - 1016
      "00000000000011100111001111000000", --  255 - 1020
      "00000000000111001110001111000000", --  256 - 1024
      "00000000000000000000000000000000", --  257 - 1028
      "00000000000000000000000000000000", --  258 - 1032
      "00010101110111000000000010001011", --  259 - 1036
      "10101100000011100000010001111000", --  260 - 1040
      "00100011110111011111111100000110", --  261 - 1044
      "00010011101000000000000000011101", --  262 - 1048
      "00100011110111011111111000001100", --  263 - 1052
      "00010011101000000000000000011011", --  264 - 1056
      "00100011110111011111110100010010", --  265 - 1060
      "00010011101000000000000000011001", --  266 - 1064
      "00100011110111101111111111111111", --  267 - 1068
      "00100011111111111111111111111111", --  268 - 1072
      "00010111110111110000000010000001", --  269 - 1076
      "00011111111000001111111101000101", --  270 - 1080
      "00010000000000000000000100001100", --  271 - 1084
      "00000000000000000000000000000000", --  272 - 1088
      "00000000000000000000000000000000", --  273 - 1092
      "00000000000000000000000000000000", --  274 - 1096
      "00000000000000000000000000000000", --  275 - 1100
      "00000000000000000000000000000000", --  276 - 1104
      "00000000000000000000000000000000", --  277 - 1108
      "00000000000000000000000000000000", --  278 - 1112
      "00000000000000000000000000000000", --  279 - 1116
      "00000000000000000000000000000000", --  280 - 1120
      "00000000000000000000000000000000", --  281 - 1124
      "00000000000000000000000000000000", --  282 - 1128
      "00000000000000000000000000000000", --  283 - 1132
      "00000000000000000000000000000000", --  284 - 1136
      "00000000000000000000000000000000", --  285 - 1140
      "00000000000000000000000000000000", --  286 - 1144
      "00000000000000000000000000000000", --  287 - 1148
      "00000000000000000000000000000000", --  288 - 1152
      "00000000000000000000000000000000", --  289 - 1156
      "00000000000000000000000000000000", --  290 - 1160
      "10001100000111010000011111100000", --  291 - 1164
      "00011111101000000000000000000011", --  292 - 1168
      "00100000000111010000000000111100", --  293 - 1172
      "00010000000000000000000000000010", --  294 - 1176
      "00100000000111010000000000000000", --  295 - 1180
      "00010100001011110000000001100110", --  296 - 1184
      "10101111101000010000011101101000", --  297 - 1188
      "10001100000111010000011111100000", --  298 - 1192
      "00011111101000000000000000000011", --  299 - 1196
      "00100000000111010000000000111100", --  300 - 1200
      "00010000000000000000000000000010", --  301 - 1204
      "00100000000111010000000000000000", --  302 - 1208
      "00010100010100000000000001011111", --  303 - 1212
      "10101111101000100000011101101100", --  304 - 1216
      "10001100000111010000011111100000", --  305 - 1220
      "00011111101000000000000000000011", --  306 - 1224
      "00100000000111010000000000111100", --  307 - 1228
      "00010000000000000000000000000010", --  308 - 1232
      "00100000000111010000000000000000", --  309 - 1236
      "00010100011100010000000001011000", --  310 - 1240
      "10101111101000110000011101110000", --  311 - 1244
      "10001100000111010000011111100000", --  312 - 1248
      "00011111101000000000000000000011", --  313 - 1252
      "00100000000111010000000000111100", --  314 - 1256
      "00010000000000000000000000000010", --  315 - 1260
      "00100000000111010000000000000000", --  316 - 1264
      "00010100100100100000000001010001", --  317 - 1268
      "10101111101001000000011101110100", --  318 - 1272
      "10001100000111010000011111100000", --  319 - 1276
      "00011111101000000000000000000011", --  320 - 1280
      "00100000000111010000000000111100", --  321 - 1284
      "00010000000000000000000000000010", --  322 - 1288
      "00100000000111010000000000000000", --  323 - 1292
      "00010100101100110000000001001010", --  324 - 1296
      "10101111101001010000011101111000", --  325 - 1300
      "10001100000111010000011111100000", --  326 - 1304
      "00011111101000000000000000000011", --  327 - 1308
      "00100000000111010000000000111100", --  328 - 1312
      "00010000000000000000000000000010", --  329 - 1316
      "00100000000111010000000000000000", --  330 - 1320
      "00010100110101000000000001000011", --  331 - 1324
      "10101111101001100000011101111100", --  332 - 1328
      "10001100000111010000011111100000", --  333 - 1332
      "00011111101000000000000000000011", --  334 - 1336
      "00100000000111010000000000111100", --  335 - 1340
      "00010000000000000000000000000010", --  336 - 1344
      "00100000000111010000000000000000", --  337 - 1348
      "00010100111101010000000000111100", --  338 - 1352
      "10101111101001110000011110000000", --  339 - 1356
      "10001100000111010000011111100000", --  340 - 1360
      "00011111101000000000000000000011", --  341 - 1364
      "00100000000111010000000000111100", --  342 - 1368
      "00010000000000000000000000000010", --  343 - 1372
      "00100000000111010000000000000000", --  344 - 1376
      "00010101000101100000000000110101", --  345 - 1380
      "10101111101010000000011110000100", --  346 - 1384
      "10001100000111010000011111100000", --  347 - 1388
      "00011111101000000000000000000011", --  348 - 1392
      "00100000000111010000000000111100", --  349 - 1396
      "00010000000000000000000000000010", --  350 - 1400
      "00100000000111010000000000000000", --  351 - 1404
      "00010101001101110000000000101110", --  352 - 1408
      "10101111101010010000011110001000", --  353 - 1412
      "10001100000111010000011111100000", --  354 - 1416
      "00011111101000000000000000000011", --  355 - 1420
      "00100000000111010000000000111100", --  356 - 1424
      "00010000000000000000000000000010", --  357 - 1428
      "00100000000111010000000000000000", --  358 - 1432
      "00010101010110000000000000100111", --  359 - 1436
      "10101111101010100000011110001100", --  360 - 1440
      "10001100000111010000011111100000", --  361 - 1444
      "00011111101000000000000000000011", --  362 - 1448
      "00100000000111010000000000111100", --  363 - 1452
      "00010000000000000000000000000010", --  364 - 1456
      "00100000000111010000000000000000", --  365 - 1460
      "00010101011110010000000000100000", --  366 - 1464
      "10101111101010110000011110010000", --  367 - 1468
      "10001100000111010000011111100000", --  368 - 1472
      "00011111101000000000000000000011", --  369 - 1476
      "00100000000111010000000000111100", --  370 - 1480
      "00010000000000000000000000000010", --  371 - 1484
      "00100000000111010000000000000000", --  372 - 1488
      "00010101100110100000000000011001", --  373 - 1492
      "10101111101011000000011110010100", --  374 - 1496
      "10001100000111010000011111100000", --  375 - 1500
      "00011111101000000000000000000011", --  376 - 1504
      "00100000000111010000000000111100", --  377 - 1508
      "00010000000000000000000000000010", --  378 - 1512
      "00100000000111010000000000000000", --  379 - 1516
      "00010101101110110000000000010010", --  380 - 1520
      "10101111101011010000011110011000", --  381 - 1524
      "10001100000111010000011111100000", --  382 - 1528
      "00011111101000000000000000000011", --  383 - 1532
      "00100000000111010000000000111100", --  384 - 1536
      "00010000000000000000000000000010", --  385 - 1540
      "00100000000111010000000000000000", --  386 - 1544
      "00010101110111000000000000001011", --  387 - 1548
      "10101111101011100000011110011100", --  388 - 1552
      "10001100000111010000011111100000", --  389 - 1556
      "00011111101000000000000000000011", --  390 - 1560
      "00100000000111010000000000111100", --  391 - 1564
      "00010000000000000000000000000010", --  392 - 1568
      "00100000000111010000000000000000", --  393 - 1572
      "00010111110111110000000000000100", --  394 - 1576
      "10101111101111100000011110100000", --  395 - 1580
      "10101100000111010000011111100000", --  396 - 1584
      "00010000000000001111111101111110", --  397 - 1588
      "10001100000111010000011111100000", --  398 - 1592
      "10001111101000010000011101101000", --  399 - 1596
      "10001100000111010000011111100000", --  400 - 1600
      "10001111101011110000011101101000", --  401 - 1604
      "00010100001011111111111111111100", --  402 - 1608
      "10001100000111010000011111100000", --  403 - 1612
      "10001111101000100000011101101100", --  404 - 1616
      "10001100000111010000011111100000", --  405 - 1620
      "10001111101100000000011101101100", --  406 - 1624
      "00010100010100001111111111111100", --  407 - 1628
      "10001100000111010000011111100000", --  408 - 1632
      "10001111101000110000011101110000", --  409 - 1636
      "10001100000111010000011111100000", --  410 - 1640
      "10001111101100010000011101110000", --  411 - 1644
      "00010100011100011111111111111100", --  412 - 1648
      "10001100000111010000011111100000", --  413 - 1652
      "10001111101001000000011101110100", --  414 - 1656
      "10001100000111010000011111100000", --  415 - 1660
      "10001111101100100000011101110100", --  416 - 1664
      "00010100100100101111111111111100", --  417 - 1668
      "10001100000111010000011111100000", --  418 - 1672
      "10001111101001010000011101111000", --  419 - 1676
      "10001100000111010000011111100000", --  420 - 1680
      "10001111101100110000011101111000", --  421 - 1684
      "00010100101100111111111111111100", --  422 - 1688
      "10001100000111010000011111100000", --  423 - 1692
      "10001111101001100000011101111100", --  424 - 1696
      "10001100000111010000011111100000", --  425 - 1700
      "10001111101101000000011101111100", --  426 - 1704
      "00010100110101001111111111111100", --  427 - 1708
      "10001100000111010000011111100000", --  428 - 1712
      "10001111101001110000011110000000", --  429 - 1716
      "10001100000111010000011111100000", --  430 - 1720
      "10001111101101010000011110000000", --  431 - 1724
      "00010100111101011111111111111100", --  432 - 1728
      "10001100000111010000011111100000", --  433 - 1732
      "10001111101010000000011110000100", --  434 - 1736
      "10001100000111010000011111100000", --  435 - 1740
      "10001111101101100000011110000100", --  436 - 1744
      "00010101000101101111111111111100", --  437 - 1748
      "10001100000111010000011111100000", --  438 - 1752
      "10001111101010010000011110001000", --  439 - 1756
      "10001100000111010000011111100000", --  440 - 1760
      "10001111101101110000011110001000", --  441 - 1764
      "00010101001101111111111111111100", --  442 - 1768
      "10001100000111010000011111100000", --  443 - 1772
      "10001111101010100000011110001100", --  444 - 1776
      "10001100000111010000011111100000", --  445 - 1780
      "10001111101110000000011110001100", --  446 - 1784
      "00010101010110001111111111111100", --  447 - 1788
      "10001100000111010000011111100000", --  448 - 1792
      "10001111101010110000011110010000", --  449 - 1796
      "10001100000111010000011111100000", --  450 - 1800
      "10001111101110010000011110010000", --  451 - 1804
      "00010101011110011111111111111100", --  452 - 1808
      "10001100000111010000011111100000", --  453 - 1812
      "10001111101011000000011110010100", --  454 - 1816
      "10001100000111010000011111100000", --  455 - 1820
      "10001111101110100000011110010100", --  456 - 1824
      "00010101100110101111111111111100", --  457 - 1828
      "10001100000111010000011111100000", --  458 - 1832
      "10001111101011010000011110011000", --  459 - 1836
      "10001100000111010000011111100000", --  460 - 1840
      "10001111101110110000011110011000", --  461 - 1844
      "00010101101110111111111111111100", --  462 - 1848
      "10001100000111010000011111100000", --  463 - 1852
      "10001111101011100000011110011100", --  464 - 1856
      "10001100000111010000011111100000", --  465 - 1860
      "10001111101111000000011110011100", --  466 - 1864
      "00010101110111001111111111111100", --  467 - 1868
      "10001100000111010000011111100000", --  468 - 1872
      "10001111101111100000011110100000", --  469 - 1876
      "10001100000111010000011111100000", --  470 - 1880
      "10001111101111110000011110100000", --  471 - 1884
      "00010111110111111111111111111100", --  472 - 1888
      "00010000000000001111111100110010", --  473 - 1892
      "00000000000000000000000000000000", --  474 - 1896
      "00000000000000000000000000000000", --  475 - 1900
      "00000000000000000000000000000000", --  476 - 1904
      "00000000000000000000000000000000", --  477 - 1908
      "00000000000000000000000000000000", --  478 - 1912
      "00000000000000000000000000000000", --  479 - 1916
      "00000000000000000000000000000000", --  480 - 1920
      "00000000000000000000000000000000", --  481 - 1924
      "00000000000000000000000000000000", --  482 - 1928
      "00000000000000000000000000000000", --  483 - 1932
      "00000000000000000000000000000000", --  484 - 1936
      "00000000000000000000000000000000", --  485 - 1940
      "00000000000000000000000000000000", --  486 - 1944
      "00000000000000000000000000000000", --  487 - 1948
      "00000000000000000000000000000000", --  488 - 1952
      "00000000000000000000000000000000", --  489 - 1956
      "00000000000000000000000000000000", --  490 - 1960
      "00000000000000000000000000000000", --  491 - 1964
      "00000000000000000000000000000000", --  492 - 1968
      "00000000000000000000000000000000", --  493 - 1972
      "00000000000000000000000000000000", --  494 - 1976
      "00000000000000000000000000000000", --  495 - 1980
      "00000000000000000000000000000000", --  496 - 1984
      "00000000000000000000000000000000", --  497 - 1988
      "00000000000000000000000000000000", --  498 - 1992
      "00000000000000000000000000000000", --  499 - 1996
      "00000000000000000000000000000000", --  500 - 2000
      "00000000000000000000000000000000", --  501 - 2004
      "00000000000000000000000000000000", --  502 - 2008
      "00000000000000000000000000000000", --  503 - 2012
      "00000000000000000000001111100111", --  504 - 2016
      "00000000000000000000000000000000", --  505 - 2020
      "00000000000000000000000000000000", --  506 - 2024
      "00000000000000000000000000000000", --  507 - 2028
      "00000000000000000000000000000000", --  508 - 2032
      "00000000000000000000000000000000", --  509 - 2036
      "00000000000000000000000000000000", --  510 - 2040
      "00000000000000000000000000000000", --  511 - 2044
      "00000000000000000000000000000000", --  512 - 2048
      "00000000000000000000000000000000", --  513 - 2052
      "00000000000000000000000000000000", --  514 - 2056
      "00000000000000000000000000000000", --  515 - 2060
      "00000000000000000000000000000000", --  516 - 2064
      "00000000000000000000000000000000", --  517 - 2068
      "00000000000000000000000000000000", --  518 - 2072
      "00000000000000000000000000000000", --  519 - 2076
      "00000000000000000000000000000000", --  520 - 2080
      "00000000000000000000000000000000", --  521 - 2084
      "00000000000000000000000000000000", --  522 - 2088
      "00000000000000000000000000000000", --  523 - 2092
      "00000000000000000000000000000000", --  524 - 2096
      "00000000000000000000000000000000", --  525 - 2100
      "00000000000000000000000000000000", --  526 - 2104
      "00000000000000000000000000000000", --  527 - 2108
      "00000000000000000000000000000000", --  528 - 2112
      "00000000000000000000000000000000", --  529 - 2116
      "00000000000000000000000000000000", --  530 - 2120
      "00000000000000000000000000000000", --  531 - 2124
      "00000000000000000000000000000000", --  532 - 2128
      "00000000000000000000000000000000", --  533 - 2132
      "00000000000000000000000000000000", --  534 - 2136
      "00000000000000000000000000000000", --  535 - 2140
      "00000000000000000000000000000000", --  536 - 2144
      "00000000000000000000000000000000", --  537 - 2148
      "00000000000000000000000000000000", --  538 - 2152
      "00000000000000000000000000000000");--  539 - 2156

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000010001001011010101";
         f_reg(4) <= "00000000001000010001000000100010";
         f_reg(5) <= "00101000001000110010100010011111";
         f_reg(6) <= "00000000001000010010000000100000";
         f_reg(7) <= "00000000000000100010100001000011";
         f_reg(8) <= "00000000101000110011000000100011";
         f_reg(9) <= "00000000010000100011100000100101";
         f_reg(10) <= "00000000000000000100000111000011";
         f_reg(11) <= "10101100000010000000010001000000";
         f_reg(12) <= "10101100000000010000010001000100";
         f_reg(13) <= "00000000100001000100100000000110";
         f_reg(14) <= "00000000111001110101000000101011";
         f_reg(15) <= "00000000110010100101100000100111";
         f_reg(16) <= "10101100000010000000010001001000";
         f_reg(17) <= "00000001000000010110000000000100";
         f_reg(18) <= "00000000000000000000000000000000";
         f_reg(19) <= "00000001100010110110100000101011";
         f_reg(20) <= "00000000000010000111000110000010";
         f_reg(21) <= "10101100000000010000010001001100";
         f_reg(22) <= "00000001001001010010100000101011";
         f_reg(23) <= "00000000001001100111100000100011";
         f_reg(24) <= "00000000100000111000000000100100";
         f_reg(25) <= "00101001110100011000100100101101";
         f_reg(26) <= "00000000100001101001000000100111";
         f_reg(27) <= "00101101000100110100100000000010";
         f_reg(28) <= "00000001101000011010000000100100";
         f_reg(29) <= "10101100000011000000010001010000";
         f_reg(30) <= "00000000000000011010100000000110";
         f_reg(31) <= "00000010010011101011000000100001";
         f_reg(32) <= "00000000101011111011100000101010";
         f_reg(33) <= "00000001011010101100000000100001";
         f_reg(34) <= "10101100000010100000010001010100";
         f_reg(35) <= "00000000000000000000000000000000";
         f_reg(36) <= "00000010011100101100100000100101";
         f_reg(37) <= "00000000000010011101010000000011";
         f_reg(38) <= "10101100000110010000010001011000";
         f_reg(39) <= "00000000110001000011000000100010";
         f_reg(40) <= "00100110111110111101010011110111";
         f_reg(41) <= "00000000101011010010100000100111";
         f_reg(42) <= "00000000000110011110010000000011";
         f_reg(43) <= "00101101011111010001011001001101";
         f_reg(44) <= "00000011011100001111000000101011";
         f_reg(45) <= "00000011000100100001000000100000";
         f_reg(46) <= "00000010100000000011100000100100";
         f_reg(47) <= "10101100000001110000010001011100";
         f_reg(48) <= "00110010101000111000000001111000";
         f_reg(49) <= "00000000010111100110000000100011";
         f_reg(50) <= "00000011010111000000100000100010";
         f_reg(51) <= "00000000110111100111000000101011";
         f_reg(52) <= "00000000010010000111100000100101";
         f_reg(53) <= "00100111001010101000000100111100";
         f_reg(54) <= "00111000101010011100000101001101";
         f_reg(55) <= "10101100000100010000010001100000";
         f_reg(56) <= "00101101110001000110110111011111";
         f_reg(57) <= "10101100000011110000010001100100";
         f_reg(58) <= "10101100000010100000010001101000";
         f_reg(59) <= "00000011110010011011100000000100";
         f_reg(60) <= "00000000011111010110100000101010";
         f_reg(61) <= "00000000001001000101100000100110";
         f_reg(62) <= "00000000110011101101100000100111";
         f_reg(63) <= "00000000000000000000000000000000";
         f_reg(64) <= "10101100000110110000010001101100";
         f_reg(65) <= "10101100000011010000010001110000";
         f_reg(66) <= "00000010111000001000000000100100";
         f_reg(67) <= "00000010011011001100000000100010";
         f_reg(68) <= "00000010110010111001000000100000";
         f_reg(69) <= "00000000000000000000000000000000";
         f_reg(70) <= "00110110000101000111000001000101";
         f_reg(71) <= "00000000000000000000000000000000";
         f_reg(72) <= "00000010100110000011100000101011";
         f_reg(73) <= "10101100000001110000010001110100";
         f_reg(74) <= "00000000000100101001001111000000";
         f_reg(75) <= "00000000000000000000000000000000";
         f_reg(76) <= "10101100000100100000010001111000";
         f_reg(77) <= "00100011111111111111111111111111";
         f_reg(78) <= "00011111111000001111111110110101";
         f_reg(79) <= "00010000000000000000000111001101";
         f_reg(80) <= "00111100000111100000001111100111";
         f_reg(81) <= "00111100000111110000001111100111";
         f_reg(82) <= "00000000000111101111010000000010";
         f_reg(83) <= "00000000000111111111110000000010";
         f_reg(84) <= "00111100000000010001001011010101";
         f_reg(85) <= "00111100000011110001001011010101";
         f_reg(86) <= "00000000001000010001000000100010";
         f_reg(87) <= "00000001111011111000000000100010";
         f_reg(88) <= "00101000001000110010100010011111";
         f_reg(89) <= "00101001111100010010100010011111";
         f_reg(90) <= "00000000001000010010000000100000";
         f_reg(91) <= "00000001111011111001000000100000";
         f_reg(92) <= "00000000000000100010100001000011";
         f_reg(93) <= "00000000000100001001100001000011";
         f_reg(94) <= "00000000101000110011000000100011";
         f_reg(95) <= "00000010011100011010000000100011";
         f_reg(96) <= "00000000010000100011100000100101";
         f_reg(97) <= "00000010000100001010100000100101";
         f_reg(98) <= "00000000000000000100000111000011";
         f_reg(99) <= "00000000000000001011000111000011";
         f_reg(100) <= "00010101000101100000000100101011";
         f_reg(101) <= "10101100000010000000010001000000";
         f_reg(102) <= "00010100001011110000000100101001";
         f_reg(103) <= "10101100000000010000010001000100";
         f_reg(104) <= "00000000100001000100100000000110";
         f_reg(105) <= "00000010010100101011100000000110";
         f_reg(106) <= "00000000111001110101000000101011";
         f_reg(107) <= "00000010101101011100000000101011";
         f_reg(108) <= "00000000110010100101100000100111";
         f_reg(109) <= "00000010100110001100100000100111";
         f_reg(110) <= "00010101000101100000000100100001";
         f_reg(111) <= "10101100000010000000010001001000";
         f_reg(112) <= "00000001000000010110000000000100";
         f_reg(113) <= "00000010110011111101000000000100";
         f_reg(114) <= "00000000000000000000000000000000";
         f_reg(115) <= "00000000000000000000000000000000";
         f_reg(116) <= "00000001100010110110100000101011";
         f_reg(117) <= "00000011010110011101100000101011";
         f_reg(118) <= "00000000000010000111000110000010";
         f_reg(119) <= "00000000000101101110000110000010";
         f_reg(120) <= "00010100001011110000000100010111";
         f_reg(121) <= "10101100000000010000010001001100";
         f_reg(122) <= "00000001001001010010100000101011";
         f_reg(123) <= "00000010111100111001100000101011";
         f_reg(124) <= "00000000001001100001000000100011";
         f_reg(125) <= "00000001111101001000000000100011";
         f_reg(126) <= "00000000100000110011100000100100";
         f_reg(127) <= "00000010010100011010100000100100";
         f_reg(128) <= "00101001110000111000100100101101";
         f_reg(129) <= "00101011100100011000100100101101";
         f_reg(130) <= "00010100011100010000000100001101";
         f_reg(131) <= "10101100000000110000010001111100";
         f_reg(132) <= "00000000100001100001100000100111";
         f_reg(133) <= "00000010010101001000100000100111";
         f_reg(134) <= "00010100011100010000000100001001";
         f_reg(135) <= "10101100000000110000010010000000";
         f_reg(136) <= "00101101000000110100100000000010";
         f_reg(137) <= "00101110110100010100100000000010";
         f_reg(138) <= "00010100011100010000000100000101";
         f_reg(139) <= "10101100000000110000010010000100";
         f_reg(140) <= "00000001101000010001100000100100";
         f_reg(141) <= "00000011011011111000100000100100";
         f_reg(142) <= "00010101100110100000000100000001";
         f_reg(143) <= "10101100000011000000010001010000";
         f_reg(144) <= "00000000000000010110000000000110";
         f_reg(145) <= "00000000000011111101000000000110";
         f_reg(146) <= "10001100000000010000010010000000";
         f_reg(147) <= "10001100000011110000010010000000";
         f_reg(148) <= "00010100001011111111111111111110";
         f_reg(149) <= "00010101000101100000000011111010";
         f_reg(150) <= "10101100000010000000010010000000";
         f_reg(151) <= "00000000001011100100000000100001";
         f_reg(152) <= "00000001111111001011000000100001";
         f_reg(153) <= "00000000101000100111000000101010";
         f_reg(154) <= "00000010011100001110000000101010";
         f_reg(155) <= "00000001011010100001000000100001";
         f_reg(156) <= "00000011001110001000000000100001";
         f_reg(157) <= "00010101010110000000000011110010";
         f_reg(158) <= "10101100000010100000010001010100";
         f_reg(159) <= "00000000000000000000000000000000";
         f_reg(160) <= "00000000000000000000000000000000";
         f_reg(161) <= "10001100000010100000010010000100";
         f_reg(162) <= "10001100000110000000010010000100";
         f_reg(163) <= "00010101010110001111111111111110";
         f_reg(164) <= "00010101000101100000000011101011";
         f_reg(165) <= "10101100000010000000010010000100";
         f_reg(166) <= "00000001010000010100000000100101";
         f_reg(167) <= "00000011000011111011000000100101";
         f_reg(168) <= "00010101010110000000000011100111";
         f_reg(169) <= "10101100000010100000010010001000";
         f_reg(170) <= "00000000000010010101010000000011";
         f_reg(171) <= "00000000000101111100010000000011";
         f_reg(172) <= "00010101000101100000000011100011";
         f_reg(173) <= "10101100000010000000010001011000";
         f_reg(174) <= "00000000110001000011000000100010";
         f_reg(175) <= "00000010100100101010000000100010";
         f_reg(176) <= "00100101110010011101010011110111";
         f_reg(177) <= "00100111100101111101010011110111";
         f_reg(178) <= "00000000101011010010100000100111";
         f_reg(179) <= "00000010011110111001100000100111";
         f_reg(180) <= "00000000000010000010010000000011";
         f_reg(181) <= "00000000000101101001010000000011";
         f_reg(182) <= "00101101011011100001011001001101";
         f_reg(183) <= "00101111001111000001011001001101";
         f_reg(184) <= "00000001001001110110100000101011";
         f_reg(185) <= "00000010111101011101100000101011";
         f_reg(186) <= "00000000010000010101100000100000";
         f_reg(187) <= "00000010000011111100100000100000";
         f_reg(188) <= "00000000011000000100100000100100";
         f_reg(189) <= "00000010001000001011100000100100";
         f_reg(190) <= "00010101001101110000000011010001";
         f_reg(191) <= "10101100000010010000010001011100";
         f_reg(192) <= "00110001100001111000000001111000";
         f_reg(193) <= "00110011010101011000000001111000";
         f_reg(194) <= "00000001011011010001000000100011";
         f_reg(195) <= "00000011001110111000000000100011";
         f_reg(196) <= "00000001010001000000100000100010";
         f_reg(197) <= "00000011000100100111100000100010";
         f_reg(198) <= "00000000110011010001100000101011";
         f_reg(199) <= "00000010100110111000100000101011";
         f_reg(200) <= "10001100000010010000010010000000";
         f_reg(201) <= "10001100000101110000010010000000";
         f_reg(202) <= "00010101001101111111111111111110";
         f_reg(203) <= "00000001011010010110000000100101";
         f_reg(204) <= "00000011001101111101000000100101";
         f_reg(205) <= "00100101000010101000000100111100";
         f_reg(206) <= "00100110110110001000000100111100";
         f_reg(207) <= "00111000101001001100000101001101";
         f_reg(208) <= "00111010011100101100000101001101";
         f_reg(209) <= "10001100000010110000010001111100";
         f_reg(210) <= "10001100000110010000010001111100";
         f_reg(211) <= "00010101011110011111111111111110";
         f_reg(212) <= "00010101011110010000000010111011";
         f_reg(213) <= "10101100000010110000010001100000";
         f_reg(214) <= "00101100011010010110110111011111";
         f_reg(215) <= "00101110001101110110110111011111";
         f_reg(216) <= "00010101100110100000000010110111";
         f_reg(217) <= "10101100000011000000010001100100";
         f_reg(218) <= "00010101010110000000000010110101";
         f_reg(219) <= "10101100000010100000010001101000";
         f_reg(220) <= "00000001101001000100000000000100";
         f_reg(221) <= "00000011011100101011000000000100";
         f_reg(222) <= "00000000111011100010100000101010";
         f_reg(223) <= "00000010101111001001100000101010";
         f_reg(224) <= "00000000001010010101100000100110";
         f_reg(225) <= "00000001111101111100100000100110";
         f_reg(226) <= "00000000110000110110000000100111";
         f_reg(227) <= "00000010100100011101000000100111";
         f_reg(228) <= "00000000000000000000000000000000";
         f_reg(229) <= "00000000000000000000000000000000";
         f_reg(230) <= "00010101100110100000000010101001";
         f_reg(231) <= "10101100000011000000010001101100";
         f_reg(232) <= "00010100101100110000000010100111";
         f_reg(233) <= "10101100000001010000010001110000";
         f_reg(234) <= "00000001000000000101000000100100";
         f_reg(235) <= "00000010110000001100000000100100";
         f_reg(236) <= "10001100000001000000010010001000";
         f_reg(237) <= "10001100000100100000010010001000";
         f_reg(238) <= "00010100100100101111111111111110";
         f_reg(239) <= "00000000100000100110100000100010";
         f_reg(240) <= "00000010010100001101100000100010";
         f_reg(241) <= "10001100000001110000010010000100";
         f_reg(242) <= "10001100000101010000010010000100";
         f_reg(243) <= "00010100111101011111111111111110";
         f_reg(244) <= "00000000111010110111000000100000";
         f_reg(245) <= "00000010101110011110000000100000";
         f_reg(246) <= "00000000000000000000000000000000";
         f_reg(247) <= "00000000000000000000000000000000";
         f_reg(248) <= "00110101010000010111000001000101";
         f_reg(249) <= "00110111000011110111000001000101";
         f_reg(250) <= "00000000000000000000000000000000";
         f_reg(251) <= "00000000000000000000000000000000";
         f_reg(252) <= "00000000001011010100100000101011";
         f_reg(253) <= "00000001111110111011100000101011";
         f_reg(254) <= "00010101001101110000000010010001";
         f_reg(255) <= "10101100000010010000010001110100";
         f_reg(256) <= "00000000000011100111001111000000";
         f_reg(257) <= "00000000000111001110001111000000";
         f_reg(258) <= "00000000000000000000000000000000";
         f_reg(259) <= "00000000000000000000000000000000";
         f_reg(260) <= "00010101110111000000000010001011";
         f_reg(261) <= "10101100000011100000010001111000";
         f_reg(262) <= "00100011110111011111111100000110";
         f_reg(263) <= "00010011101000000000000000011101";
         f_reg(264) <= "00100011110111011111111000001100";
         f_reg(265) <= "00010011101000000000000000011011";
         f_reg(266) <= "00100011110111011111110100010010";
         f_reg(267) <= "00010011101000000000000000011001";
         f_reg(268) <= "00100011110111101111111111111111";
         f_reg(269) <= "00100011111111111111111111111111";
         f_reg(270) <= "00010111110111110000000010000001";
         f_reg(271) <= "00011111111000001111111101000101";
         f_reg(272) <= "00010000000000000000000100001100";
         f_reg(273) <= "00000000000000000000000000000000";
         f_reg(274) <= "00000000000000000000000000000000";
         f_reg(275) <= "00000000000000000000000000000000";
         f_reg(276) <= "00000000000000000000000000000000";
         f_reg(277) <= "00000000000000000000000000000000";
         f_reg(278) <= "00000000000000000000000000000000";
         f_reg(279) <= "00000000000000000000000000000000";
         f_reg(280) <= "00000000000000000000000000000000";
         f_reg(281) <= "00000000000000000000000000000000";
         f_reg(282) <= "00000000000000000000000000000000";
         f_reg(283) <= "00000000000000000000000000000000";
         f_reg(284) <= "00000000000000000000000000000000";
         f_reg(285) <= "00000000000000000000000000000000";
         f_reg(286) <= "00000000000000000000000000000000";
         f_reg(287) <= "00000000000000000000000000000000";
         f_reg(288) <= "00000000000000000000000000000000";
         f_reg(289) <= "00000000000000000000000000000000";
         f_reg(290) <= "00000000000000000000000000000000";
         f_reg(291) <= "00000000000000000000000000000000";
         f_reg(292) <= "10001100000111010000011111100000";
         f_reg(293) <= "00011111101000000000000000000011";
         f_reg(294) <= "00100000000111010000000000111100";
         f_reg(295) <= "00010000000000000000000000000010";
         f_reg(296) <= "00100000000111010000000000000000";
         f_reg(297) <= "00010100001011110000000001100110";
         f_reg(298) <= "10101111101000010000011101101000";
         f_reg(299) <= "10001100000111010000011111100000";
         f_reg(300) <= "00011111101000000000000000000011";
         f_reg(301) <= "00100000000111010000000000111100";
         f_reg(302) <= "00010000000000000000000000000010";
         f_reg(303) <= "00100000000111010000000000000000";
         f_reg(304) <= "00010100010100000000000001011111";
         f_reg(305) <= "10101111101000100000011101101100";
         f_reg(306) <= "10001100000111010000011111100000";
         f_reg(307) <= "00011111101000000000000000000011";
         f_reg(308) <= "00100000000111010000000000111100";
         f_reg(309) <= "00010000000000000000000000000010";
         f_reg(310) <= "00100000000111010000000000000000";
         f_reg(311) <= "00010100011100010000000001011000";
         f_reg(312) <= "10101111101000110000011101110000";
         f_reg(313) <= "10001100000111010000011111100000";
         f_reg(314) <= "00011111101000000000000000000011";
         f_reg(315) <= "00100000000111010000000000111100";
         f_reg(316) <= "00010000000000000000000000000010";
         f_reg(317) <= "00100000000111010000000000000000";
         f_reg(318) <= "00010100100100100000000001010001";
         f_reg(319) <= "10101111101001000000011101110100";
         f_reg(320) <= "10001100000111010000011111100000";
         f_reg(321) <= "00011111101000000000000000000011";
         f_reg(322) <= "00100000000111010000000000111100";
         f_reg(323) <= "00010000000000000000000000000010";
         f_reg(324) <= "00100000000111010000000000000000";
         f_reg(325) <= "00010100101100110000000001001010";
         f_reg(326) <= "10101111101001010000011101111000";
         f_reg(327) <= "10001100000111010000011111100000";
         f_reg(328) <= "00011111101000000000000000000011";
         f_reg(329) <= "00100000000111010000000000111100";
         f_reg(330) <= "00010000000000000000000000000010";
         f_reg(331) <= "00100000000111010000000000000000";
         f_reg(332) <= "00010100110101000000000001000011";
         f_reg(333) <= "10101111101001100000011101111100";
         f_reg(334) <= "10001100000111010000011111100000";
         f_reg(335) <= "00011111101000000000000000000011";
         f_reg(336) <= "00100000000111010000000000111100";
         f_reg(337) <= "00010000000000000000000000000010";
         f_reg(338) <= "00100000000111010000000000000000";
         f_reg(339) <= "00010100111101010000000000111100";
         f_reg(340) <= "10101111101001110000011110000000";
         f_reg(341) <= "10001100000111010000011111100000";
         f_reg(342) <= "00011111101000000000000000000011";
         f_reg(343) <= "00100000000111010000000000111100";
         f_reg(344) <= "00010000000000000000000000000010";
         f_reg(345) <= "00100000000111010000000000000000";
         f_reg(346) <= "00010101000101100000000000110101";
         f_reg(347) <= "10101111101010000000011110000100";
         f_reg(348) <= "10001100000111010000011111100000";
         f_reg(349) <= "00011111101000000000000000000011";
         f_reg(350) <= "00100000000111010000000000111100";
         f_reg(351) <= "00010000000000000000000000000010";
         f_reg(352) <= "00100000000111010000000000000000";
         f_reg(353) <= "00010101001101110000000000101110";
         f_reg(354) <= "10101111101010010000011110001000";
         f_reg(355) <= "10001100000111010000011111100000";
         f_reg(356) <= "00011111101000000000000000000011";
         f_reg(357) <= "00100000000111010000000000111100";
         f_reg(358) <= "00010000000000000000000000000010";
         f_reg(359) <= "00100000000111010000000000000000";
         f_reg(360) <= "00010101010110000000000000100111";
         f_reg(361) <= "10101111101010100000011110001100";
         f_reg(362) <= "10001100000111010000011111100000";
         f_reg(363) <= "00011111101000000000000000000011";
         f_reg(364) <= "00100000000111010000000000111100";
         f_reg(365) <= "00010000000000000000000000000010";
         f_reg(366) <= "00100000000111010000000000000000";
         f_reg(367) <= "00010101011110010000000000100000";
         f_reg(368) <= "10101111101010110000011110010000";
         f_reg(369) <= "10001100000111010000011111100000";
         f_reg(370) <= "00011111101000000000000000000011";
         f_reg(371) <= "00100000000111010000000000111100";
         f_reg(372) <= "00010000000000000000000000000010";
         f_reg(373) <= "00100000000111010000000000000000";
         f_reg(374) <= "00010101100110100000000000011001";
         f_reg(375) <= "10101111101011000000011110010100";
         f_reg(376) <= "10001100000111010000011111100000";
         f_reg(377) <= "00011111101000000000000000000011";
         f_reg(378) <= "00100000000111010000000000111100";
         f_reg(379) <= "00010000000000000000000000000010";
         f_reg(380) <= "00100000000111010000000000000000";
         f_reg(381) <= "00010101101110110000000000010010";
         f_reg(382) <= "10101111101011010000011110011000";
         f_reg(383) <= "10001100000111010000011111100000";
         f_reg(384) <= "00011111101000000000000000000011";
         f_reg(385) <= "00100000000111010000000000111100";
         f_reg(386) <= "00010000000000000000000000000010";
         f_reg(387) <= "00100000000111010000000000000000";
         f_reg(388) <= "00010101110111000000000000001011";
         f_reg(389) <= "10101111101011100000011110011100";
         f_reg(390) <= "10001100000111010000011111100000";
         f_reg(391) <= "00011111101000000000000000000011";
         f_reg(392) <= "00100000000111010000000000111100";
         f_reg(393) <= "00010000000000000000000000000010";
         f_reg(394) <= "00100000000111010000000000000000";
         f_reg(395) <= "00010111110111110000000000000100";
         f_reg(396) <= "10101111101111100000011110100000";
         f_reg(397) <= "10101100000111010000011111100000";
         f_reg(398) <= "00010000000000001111111101111110";
         f_reg(399) <= "10001100000111010000011111100000";
         f_reg(400) <= "10001111101000010000011101101000";
         f_reg(401) <= "10001100000111010000011111100000";
         f_reg(402) <= "10001111101011110000011101101000";
         f_reg(403) <= "00010100001011111111111111111100";
         f_reg(404) <= "10001100000111010000011111100000";
         f_reg(405) <= "10001111101000100000011101101100";
         f_reg(406) <= "10001100000111010000011111100000";
         f_reg(407) <= "10001111101100000000011101101100";
         f_reg(408) <= "00010100010100001111111111111100";
         f_reg(409) <= "10001100000111010000011111100000";
         f_reg(410) <= "10001111101000110000011101110000";
         f_reg(411) <= "10001100000111010000011111100000";
         f_reg(412) <= "10001111101100010000011101110000";
         f_reg(413) <= "00010100011100011111111111111100";
         f_reg(414) <= "10001100000111010000011111100000";
         f_reg(415) <= "10001111101001000000011101110100";
         f_reg(416) <= "10001100000111010000011111100000";
         f_reg(417) <= "10001111101100100000011101110100";
         f_reg(418) <= "00010100100100101111111111111100";
         f_reg(419) <= "10001100000111010000011111100000";
         f_reg(420) <= "10001111101001010000011101111000";
         f_reg(421) <= "10001100000111010000011111100000";
         f_reg(422) <= "10001111101100110000011101111000";
         f_reg(423) <= "00010100101100111111111111111100";
         f_reg(424) <= "10001100000111010000011111100000";
         f_reg(425) <= "10001111101001100000011101111100";
         f_reg(426) <= "10001100000111010000011111100000";
         f_reg(427) <= "10001111101101000000011101111100";
         f_reg(428) <= "00010100110101001111111111111100";
         f_reg(429) <= "10001100000111010000011111100000";
         f_reg(430) <= "10001111101001110000011110000000";
         f_reg(431) <= "10001100000111010000011111100000";
         f_reg(432) <= "10001111101101010000011110000000";
         f_reg(433) <= "00010100111101011111111111111100";
         f_reg(434) <= "10001100000111010000011111100000";
         f_reg(435) <= "10001111101010000000011110000100";
         f_reg(436) <= "10001100000111010000011111100000";
         f_reg(437) <= "10001111101101100000011110000100";
         f_reg(438) <= "00010101000101101111111111111100";
         f_reg(439) <= "10001100000111010000011111100000";
         f_reg(440) <= "10001111101010010000011110001000";
         f_reg(441) <= "10001100000111010000011111100000";
         f_reg(442) <= "10001111101101110000011110001000";
         f_reg(443) <= "00010101001101111111111111111100";
         f_reg(444) <= "10001100000111010000011111100000";
         f_reg(445) <= "10001111101010100000011110001100";
         f_reg(446) <= "10001100000111010000011111100000";
         f_reg(447) <= "10001111101110000000011110001100";
         f_reg(448) <= "00010101010110001111111111111100";
         f_reg(449) <= "10001100000111010000011111100000";
         f_reg(450) <= "10001111101010110000011110010000";
         f_reg(451) <= "10001100000111010000011111100000";
         f_reg(452) <= "10001111101110010000011110010000";
         f_reg(453) <= "00010101011110011111111111111100";
         f_reg(454) <= "10001100000111010000011111100000";
         f_reg(455) <= "10001111101011000000011110010100";
         f_reg(456) <= "10001100000111010000011111100000";
         f_reg(457) <= "10001111101110100000011110010100";
         f_reg(458) <= "00010101100110101111111111111100";
         f_reg(459) <= "10001100000111010000011111100000";
         f_reg(460) <= "10001111101011010000011110011000";
         f_reg(461) <= "10001100000111010000011111100000";
         f_reg(462) <= "10001111101110110000011110011000";
         f_reg(463) <= "00010101101110111111111111111100";
         f_reg(464) <= "10001100000111010000011111100000";
         f_reg(465) <= "10001111101011100000011110011100";
         f_reg(466) <= "10001100000111010000011111100000";
         f_reg(467) <= "10001111101111000000011110011100";
         f_reg(468) <= "00010101110111001111111111111100";
         f_reg(469) <= "10001100000111010000011111100000";
         f_reg(470) <= "10001111101111100000011110100000";
         f_reg(471) <= "10001100000111010000011111100000";
         f_reg(472) <= "10001111101111110000011110100000";
         f_reg(473) <= "00010111110111111111111111111100";
         f_reg(474) <= "00010000000000001111111100110010";
         f_reg(475) <= "00000000000000000000000000000000";
         f_reg(476) <= "00000000000000000000000000000000";
         f_reg(477) <= "00000000000000000000000000000000";
         f_reg(478) <= "00000000000000000000000000000000";
         f_reg(479) <= "00000000000000000000000000000000";
         f_reg(480) <= "00000000000000000000000000000000";
         f_reg(481) <= "00000000000000000000000000000000";
         f_reg(482) <= "00000000000000000000000000000000";
         f_reg(483) <= "00000000000000000000000000000000";
         f_reg(484) <= "00000000000000000000000000000000";
         f_reg(485) <= "00000000000000000000000000000000";
         f_reg(486) <= "00000000000000000000000000000000";
         f_reg(487) <= "00000000000000000000000000000000";
         f_reg(488) <= "00000000000000000000000000000000";
         f_reg(489) <= "00000000000000000000000000000000";
         f_reg(490) <= "00000000000000000000000000000000";
         f_reg(491) <= "00000000000000000000000000000000";
         f_reg(492) <= "00000000000000000000000000000000";
         f_reg(493) <= "00000000000000000000000000000000";
         f_reg(494) <= "00000000000000000000000000000000";
         f_reg(495) <= "00000000000000000000000000000000";
         f_reg(496) <= "00000000000000000000000000000000";
         f_reg(497) <= "00000000000000000000000000000000";
         f_reg(498) <= "00000000000000000000000000000000";
         f_reg(499) <= "00000000000000000000000000000000";
         f_reg(500) <= "00000000000000000000000000000000";
         f_reg(501) <= "00000000000000000000000000000000";
         f_reg(502) <= "00000000000000000000000000000000";
         f_reg(503) <= "00000000000000000000000000000000";
         f_reg(504) <= "00000000000000000000000000000000";
         f_reg(505) <= "00000000000000000000001111100111";
         f_reg(506) <= "00000000000000000000000000000000";
         f_reg(507) <= "00000000000000000000000000000000";
         f_reg(508) <= "00000000000000000000000000000000";
         f_reg(509) <= "00000000000000000000000000000000";
         f_reg(510) <= "00000000000000000000000000000000";
         f_reg(511) <= "00000000000000000000000000000000";
         f_reg(512) <= "00000000000000000000000000000000";
         f_reg(513) <= "00000000000000000000000000000000";
         f_reg(514) <= "00000000000000000000000000000000";
         f_reg(515) <= "00000000000000000000000000000000";
         f_reg(516) <= "00000000000000000000000000000000";
         f_reg(517) <= "00000000000000000000000000000000";
         f_reg(518) <= "00000000000000000000000000000000";
         f_reg(519) <= "00000000000000000000000000000000";
         f_reg(520) <= "00000000000000000000000000000000";
         f_reg(521) <= "00000000000000000000000000000000";
         f_reg(522) <= "00000000000000000000000000000000";
         f_reg(523) <= "00000000000000000000000000000000";
         f_reg(524) <= "00000000000000000000000000000000";
         f_reg(525) <= "00000000000000000000000000000000";
         f_reg(526) <= "00000000000000000000000000000000";
         f_reg(527) <= "00000000000000000000000000000000";
         f_reg(528) <= "00000000000000000000000000000000";
         f_reg(529) <= "00000000000000000000000000000000";
         f_reg(530) <= "00000000000000000000000000000000";
         f_reg(531) <= "00000000000000000000000000000000";
         f_reg(532) <= "00000000000000000000000000000000";
         f_reg(533) <= "00000000000000000000000000000000";
         f_reg(534) <= "00000000000000000000000000000000";
         f_reg(535) <= "00000000000000000000000000000000";
         f_reg(536) <= "00000000000000000000000000000000";
         f_reg(537) <= "00000000000000000000000000000000";
         f_reg(538) <= "00000000000000000000000000000000";
         f_reg(539) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 4821
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SUB R2 R1 R1
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SLTI R3 R1 10399
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- ADD R4 R1 R1
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SRA R5 R2 1
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- SUBU R6 R5 R3
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- OR R7 R2 R2
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- SRA R8 R0 7
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- SW R8 R0 1088
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- SW R1 R0 1092
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- SRLV R9 R4 R4
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- SLTU R10 R7 R7
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- NOR R11 R6 R10
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- SW R8 R0 1096
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- SLLV R12 R1 R8
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- NOP
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SLTU R13 R12 R11
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- SRL R14 R8 6
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SW R1 R0 1100
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- SLTU R5 R9 R5
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- SUBU R15 R1 R6
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- AND R16 R4 R3
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- SLTI R17 R14 -30419
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- NOR R18 R4 R6
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- SLTIU R19 R8 18434
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- AND R20 R13 R1
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- SW R12 R0 1104
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- SRLV R21 R1 R0
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- ADDU R22 R18 R14
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- SLT R23 R5 R15
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- ADDU R24 R11 R10
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- SW R10 R0 1108
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- NOP
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- OR R25 R19 R18
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- SRA R26 R9 16
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- SW R25 R0 1112
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- SUB R6 R6 R4
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- ADDIU R27 R23 -11017
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- NOR R5 R5 R13
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- SRA R28 R25 16
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SLTIU R29 R11 5709
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- SLTU R30 R27 R16
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- ADD R2 R24 R18
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- AND R7 R20 R0
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- SW R7 R0 1116
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- ANDI R3 R21 -32648
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- SUBU R12 R2 R30
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- SUB R1 R26 R28
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SLTU R14 R6 R30
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- OR R15 R2 R8
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- ADDIU R10 R25 -32452
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- XORI R9 R5 -16051
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SW R17 R0 1120
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- SLTIU R4 R14 28127
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SW R15 R0 1124
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- SW R10 R0 1128
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- SLLV R23 R9 R30
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SLT R13 R3 R29
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- XOR R11 R1 R4
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- NOR R27 R6 R14
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- NOP
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- SW R27 R0 1132
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- SW R13 R0 1136
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- AND R16 R23 R0
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- SUB R24 R19 R12
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- ADD R18 R22 R11
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- NOP
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- ORI R20 R16 28741
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- NOP
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- SLTU R7 R20 R24
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SW R7 R0 1140
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- SLL R18 R18 15
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- NOP
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- SW R18 R0 1144
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- BGTZ R31 -75
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- BEQ R0 R0 461
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- LUI R30 999
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- LUI R31 999
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- LUI R1 4821
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- LUI R15 4821
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- SUB R2 R1 R1
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SUB R16 R15 R15
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- SLTI R3 R1 10399
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- SLTI R17 R15 10399
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- ADD R4 R1 R1
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- ADD R18 R15 R15
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- SRA R5 R2 1
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- SRA R19 R16 1
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- SUBU R6 R5 R3
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- SUBU R20 R19 R17
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- OR R7 R2 R2
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- OR R21 R16 R16
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SRA R8 R0 7
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- SRA R22 R0 7
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- BNE R8 R22 299
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- SW R8 R0 1088
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- BNE R1 R15 297
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SW R1 R0 1092
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- SRLV R9 R4 R4
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- SRLV R23 R18 R18
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- SLTU R10 R7 R7
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- SLTU R24 R21 R21
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- NOR R11 R6 R10
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- NOR R25 R20 R24
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- BNE R8 R22 289
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- SW R8 R0 1096
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- SLLV R12 R1 R8
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- SLLV R26 R15 R22
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- NOP
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- NOP
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- SLTU R13 R12 R11
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- SLTU R27 R26 R25
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- SRL R14 R8 6
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- SRL R28 R22 6
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- BNE R1 R15 279
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- SW R1 R0 1100
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- SLTU R5 R9 R5
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- SLTU R19 R23 R19
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SUBU R2 R1 R6
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- SUBU R16 R15 R20
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- AND R7 R4 R3
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- AND R21 R18 R17
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SLTI R3 R14 -30419
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- SLTI R17 R28 -30419
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- BNE R3 R17 269
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- SW R3 R0 1148
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- NOR R3 R4 R6
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- NOR R17 R18 R20
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- BNE R3 R17 265
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- SW R3 R0 1152
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- SLTIU R3 R8 18434
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- SLTIU R17 R22 18434
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- BNE R3 R17 261
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- SW R3 R0 1156
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- AND R3 R13 R1
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- AND R17 R27 R15
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- BNE R12 R26 257
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- SW R12 R0 1104
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- SRLV R12 R1 R0
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- SRLV R26 R15 R0
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- LW R1 R0 1152
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- LW R15 R0 1152
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- BNE R1 R15 -2
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- BNE R8 R22 250
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- SW R8 R0 1152
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- ADDU R8 R1 R14
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- ADDU R22 R15 R28
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- SLT R14 R5 R2
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- SLT R28 R19 R16
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- ADDU R2 R11 R10
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- ADDU R16 R25 R24
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- BNE R10 R24 242
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- SW R10 R0 1108
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- NOP
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- NOP
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- LW R10 R0 1156
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- LW R24 R0 1156
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- BNE R10 R24 -2
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- BNE R8 R22 235
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- SW R8 R0 1156
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- OR R8 R10 R1
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- OR R22 R24 R15
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- BNE R10 R24 231
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- SW R10 R0 1160
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- SRA R10 R9 16
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- SRA R24 R23 16
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- BNE R8 R22 227
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- SW R8 R0 1112
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- SUB R6 R6 R4
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- SUB R20 R20 R18
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- ADDIU R9 R14 -11017
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- ADDIU R23 R28 -11017
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- NOR R5 R5 R13
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- NOR R19 R19 R27
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- SRA R4 R8 16
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- SRA R18 R22 16
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SLTIU R14 R11 5709
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- SLTIU R28 R25 5709
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- SLTU R13 R9 R7
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- SLTU R27 R23 R21
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- ADD R11 R2 R1
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- ADD R25 R16 R15
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- AND R9 R3 R0
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- AND R23 R17 R0
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- BNE R9 R23 209
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- SW R9 R0 1116
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- ANDI R7 R12 -32648
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- ANDI R21 R26 -32648
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- SUBU R2 R11 R13
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- SUBU R16 R25 R27
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- SUB R1 R10 R4
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- SUB R15 R24 R18
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- SLTU R3 R6 R13
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- SLTU R17 R20 R27
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- LW R9 R0 1152
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- LW R23 R0 1152
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- BNE R9 R23 -2
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- OR R12 R11 R9
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- OR R26 R25 R23
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- ADDIU R10 R8 -32452
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- ADDIU R24 R22 -32452
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- XORI R4 R5 -16051
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- XORI R18 R19 -16051
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- LW R11 R0 1148
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- LW R25 R0 1148
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- BNE R11 R25 -2
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- BNE R11 R25 187
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- SW R11 R0 1120
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- SLTIU R9 R3 28127
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- SLTIU R23 R17 28127
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- BNE R12 R26 183
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- SW R12 R0 1124
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- BNE R10 R24 181
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- SW R10 R0 1128
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- SLLV R8 R4 R13
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- SLLV R22 R18 R27
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- SLT R5 R7 R14
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- SLT R19 R21 R28
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- XOR R11 R1 R9
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- XOR R25 R15 R23
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- NOR R12 R6 R3
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- NOR R26 R20 R17
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- NOP
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- NOP
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- BNE R12 R26 169
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- SW R12 R0 1132
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- BNE R5 R19 167
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- SW R5 R0 1136
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- AND R10 R8 R0
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- AND R24 R22 R0
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- LW R4 R0 1160
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- LW R18 R0 1160
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- BNE R4 R18 -2
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- SUB R13 R4 R2
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- SUB R27 R18 R16
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- LW R7 R0 1156
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- LW R21 R0 1156
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- BNE R7 R21 -2
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- ADD R14 R7 R11
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- ADD R28 R21 R25
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- NOP
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- NOP
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- ORI R1 R10 28741
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- ORI R15 R24 28741
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- NOP
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- NOP
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- SLTU R9 R1 R13
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- SLTU R23 R15 R27
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- BNE R9 R23 145
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- SW R9 R0 1140
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- SLL R14 R14 15
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- SLL R28 R28 15
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- NOP
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- NOP
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- BNE R14 R28 139
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- SW R14 R0 1144
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- BEQ R29 R0 29
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- BEQ R29 R0 27
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- BEQ R29 R0 25
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- BNE R30 R31 129
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- BGTZ R31 -187
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- BEQ R0 R0 268
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- NOP
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- NOP
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- NOP
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- NOP
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- NOP
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- NOP
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- NOP
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- NOP
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- NOP
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- NOP
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- NOP
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- NOP
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- NOP
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- NOP
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- NOP
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- NOP
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- NOP
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- NOP
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- NOP
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- SW R1 R29 1896
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- SW R2 R29 1900
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- SW R3 R29 1904
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- SW R4 R29 1908
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- SW R5 R29 1912
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- SW R6 R29 1916
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- SW R7 R29 1920
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- SW R8 R29 1924
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- SW R9 R29 1928
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- SW R10 R29 1932
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- SW R11 R29 1936
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- SW R12 R29 1940
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- SW R13 R29 1944
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- SW R14 R29 1948
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- SW R30 R29 1952
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- SW R29 R0 2016
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- BEQ R0 R0 -130
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- LW R1 R29 1896
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- LW R15 R29 1896
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- LW R2 R29 1900
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- LW R16 R29 1900
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- LW R3 R29 1904
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- LW R17 R29 1904
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- LW R4 R29 1908
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- LW R18 R29 1908
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- LW R5 R29 1912
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- LW R19 R29 1912
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R6 R29 1916
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- LW R20 R29 1916
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- LW R7 R29 1920
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- LW R21 R29 1920
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- LW R8 R29 1924
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- LW R22 R29 1924
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- LW R9 R29 1928
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- LW R23 R29 1928
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- LW R10 R29 1932
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- LW R24 R29 1932
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- LW R11 R29 1936
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- LW R25 R29 1936
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- LW R12 R29 1940
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- LW R26 R29 1940
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- LW R13 R29 1944
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- LW R27 R29 1944
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- LW R14 R29 1948
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- LW R28 R29 1948
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- LW R30 R29 1952
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- LW R29 R0 2016
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- LW R31 R29 1952
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- BEQ R0 R0 -206
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- NOP
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- NOP
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- NOP
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- NOP
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- NOP
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- NOP
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- NOP
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- NOP
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- NOP
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- NOP
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- NOP
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- NOP
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- NOP
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- NOP
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- NOP
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- NOP
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- NOP
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- NOP
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- NOP
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- NOP
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- NOP
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- NOP
                        f_data <= f_reg(496);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(497) =>
                        -- NOP
                        f_data <= f_reg(497);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(498) =>
                        -- NOP
                        f_data <= f_reg(498);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(499) =>
                        -- NOP
                        f_data <= f_reg(499);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(500) =>
                        -- NOP
                        f_data <= f_reg(500);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(501) =>
                        -- NOP
                        f_data <= f_reg(501);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(502) =>
                        -- NOP
                        f_data <= f_reg(502);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(503) =>
                        -- NOP
                        f_data <= f_reg(503);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(504) =>
                        -- NOP
                        f_data <= f_reg(504);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(505) =>
                        -- NOP
                        f_data <= f_reg(505);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(506) =>
                        -- NOP
                        f_data <= f_reg(506);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(507) =>
                        -- NOP
                        f_data <= f_reg(507);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(508) =>
                        -- NOP
                        f_data <= f_reg(508);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(509) =>
                        -- NOP
                        f_data <= f_reg(509);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(510) =>
                        -- NOP
                        f_data <= f_reg(510);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(511) =>
                        -- NOP
                        f_data <= f_reg(511);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(512) =>
                        -- NOP
                        f_data <= f_reg(512);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(513) =>
                        -- NOP
                        f_data <= f_reg(513);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(514) =>
                        -- NOP
                        f_data <= f_reg(514);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(515) =>
                        -- NOP
                        f_data <= f_reg(515);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(516) =>
                        -- NOP
                        f_data <= f_reg(516);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(517) =>
                        -- NOP
                        f_data <= f_reg(517);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(518) =>
                        -- NOP
                        f_data <= f_reg(518);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(519) =>
                        -- NOP
                        f_data <= f_reg(519);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(520) =>
                        -- NOP
                        f_data <= f_reg(520);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(521) =>
                        -- NOP
                        f_data <= f_reg(521);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(522) =>
                        -- NOP
                        f_data <= f_reg(522);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(523) =>
                        -- NOP
                        f_data <= f_reg(523);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(524) =>
                        -- NOP
                        f_data <= f_reg(524);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(525) =>
                        -- NOP
                        f_data <= f_reg(525);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(526) =>
                        -- NOP
                        f_data <= f_reg(526);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(527) =>
                        -- NOP
                        f_data <= f_reg(527);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(528) =>
                        -- NOP
                        f_data <= f_reg(528);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(529) =>
                        -- NOP
                        f_data <= f_reg(529);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(530) =>
                        -- NOP
                        f_data <= f_reg(530);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(531) =>
                        -- NOP
                        f_data <= f_reg(531);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(532) =>
                        -- NOP
                        f_data <= f_reg(532);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(533) =>
                        -- NOP
                        f_data <= f_reg(533);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(534) =>
                        -- NOP
                        f_data <= f_reg(534);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(535) =>
                        -- NOP
                        f_data <= f_reg(535);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(536) =>
                        -- NOP
                        f_data <= f_reg(536);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(537) =>
                        -- NOP
                        f_data <= f_reg(537);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(538) =>
                        -- NOP
                        f_data <= f_reg(538);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(539) =>
                        -- NOP
                        f_data <= f_reg(539);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(540) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010001001011010101";
                        f_reg(4) <= "00000000001000010001000000100010";
                        f_reg(5) <= "00101000001000110010100010011111";
                        f_reg(6) <= "00000000001000010010000000100000";
                        f_reg(7) <= "00000000000000100010100001000011";
                        f_reg(8) <= "00000000101000110011000000100011";
                        f_reg(9) <= "00000000010000100011100000100101";
                        f_reg(10) <= "00000000000000000100000111000011";
                        f_reg(11) <= "10101100000010000000010001000000";
                        f_reg(12) <= "10101100000000010000010001000100";
                        f_reg(13) <= "00000000100001000100100000000110";
                        f_reg(14) <= "00000000111001110101000000101011";
                        f_reg(15) <= "00000000110010100101100000100111";
                        f_reg(16) <= "10101100000010000000010001001000";
                        f_reg(17) <= "00000001000000010110000000000100";
                        f_reg(18) <= "00000000000000000000000000000000";
                        f_reg(19) <= "00000001100010110110100000101011";
                        f_reg(20) <= "00000000000010000111000110000010";
                        f_reg(21) <= "10101100000000010000010001001100";
                        f_reg(22) <= "00000001001001010010100000101011";
                        f_reg(23) <= "00000000001001100111100000100011";
                        f_reg(24) <= "00000000100000111000000000100100";
                        f_reg(25) <= "00101001110100011000100100101101";
                        f_reg(26) <= "00000000100001101001000000100111";
                        f_reg(27) <= "00101101000100110100100000000010";
                        f_reg(28) <= "00000001101000011010000000100100";
                        f_reg(29) <= "10101100000011000000010001010000";
                        f_reg(30) <= "00000000000000011010100000000110";
                        f_reg(31) <= "00000010010011101011000000100001";
                        f_reg(32) <= "00000000101011111011100000101010";
                        f_reg(33) <= "00000001011010101100000000100001";
                        f_reg(34) <= "10101100000010100000010001010100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000010011100101100100000100101";
                        f_reg(37) <= "00000000000010011101010000000011";
                        f_reg(38) <= "10101100000110010000010001011000";
                        f_reg(39) <= "00000000110001000011000000100010";
                        f_reg(40) <= "00100110111110111101010011110111";
                        f_reg(41) <= "00000000101011010010100000100111";
                        f_reg(42) <= "00000000000110011110010000000011";
                        f_reg(43) <= "00101101011111010001011001001101";
                        f_reg(44) <= "00000011011100001111000000101011";
                        f_reg(45) <= "00000011000100100001000000100000";
                        f_reg(46) <= "00000010100000000011100000100100";
                        f_reg(47) <= "10101100000001110000010001011100";
                        f_reg(48) <= "00110010101000111000000001111000";
                        f_reg(49) <= "00000000010111100110000000100011";
                        f_reg(50) <= "00000011010111000000100000100010";
                        f_reg(51) <= "00000000110111100111000000101011";
                        f_reg(52) <= "00000000010010000111100000100101";
                        f_reg(53) <= "00100111001010101000000100111100";
                        f_reg(54) <= "00111000101010011100000101001101";
                        f_reg(55) <= "10101100000100010000010001100000";
                        f_reg(56) <= "00101101110001000110110111011111";
                        f_reg(57) <= "10101100000011110000010001100100";
                        f_reg(58) <= "10101100000010100000010001101000";
                        f_reg(59) <= "00000011110010011011100000000100";
                        f_reg(60) <= "00000000011111010110100000101010";
                        f_reg(61) <= "00000000001001000101100000100110";
                        f_reg(62) <= "00000000110011101101100000100111";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000110110000010001101100";
                        f_reg(65) <= "10101100000011010000010001110000";
                        f_reg(66) <= "00000010111000001000000000100100";
                        f_reg(67) <= "00000010011011001100000000100010";
                        f_reg(68) <= "00000010110010111001000000100000";
                        f_reg(69) <= "00000000000000000000000000000000";
                        f_reg(70) <= "00110110000101000111000001000101";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000010100110000011100000101011";
                        f_reg(73) <= "10101100000001110000010001110100";
                        f_reg(74) <= "00000000000100101001001111000000";
                        f_reg(75) <= "00000000000000000000000000000000";
                        f_reg(76) <= "10101100000100100000010001111000";
                        f_reg(77) <= "00100011111111111111111111111111";
                        f_reg(78) <= "00011111111000001111111110110101";
                        f_reg(79) <= "00010000000000000000000111001101";
                        f_reg(80) <= "00111100000111100000001111100111";
                        f_reg(81) <= "00111100000111110000001111100111";
                        f_reg(82) <= "00000000000111101111010000000010";
                        f_reg(83) <= "00000000000111111111110000000010";
                        f_reg(84) <= "00111100000000010001001011010101";
                        f_reg(85) <= "00111100000011110001001011010101";
                        f_reg(86) <= "00000000001000010001000000100010";
                        f_reg(87) <= "00000001111011111000000000100010";
                        f_reg(88) <= "00101000001000110010100010011111";
                        f_reg(89) <= "00101001111100010010100010011111";
                        f_reg(90) <= "00000000001000010010000000100000";
                        f_reg(91) <= "00000001111011111001000000100000";
                        f_reg(92) <= "00000000000000100010100001000011";
                        f_reg(93) <= "00000000000100001001100001000011";
                        f_reg(94) <= "00000000101000110011000000100011";
                        f_reg(95) <= "00000010011100011010000000100011";
                        f_reg(96) <= "00000000010000100011100000100101";
                        f_reg(97) <= "00000010000100001010100000100101";
                        f_reg(98) <= "00000000000000000100000111000011";
                        f_reg(99) <= "00000000000000001011000111000011";
                        f_reg(100) <= "00010101000101100000000100101011";
                        f_reg(101) <= "10101100000010000000010001000000";
                        f_reg(102) <= "00010100001011110000000100101001";
                        f_reg(103) <= "10101100000000010000010001000100";
                        f_reg(104) <= "00000000100001000100100000000110";
                        f_reg(105) <= "00000010010100101011100000000110";
                        f_reg(106) <= "00000000111001110101000000101011";
                        f_reg(107) <= "00000010101101011100000000101011";
                        f_reg(108) <= "00000000110010100101100000100111";
                        f_reg(109) <= "00000010100110001100100000100111";
                        f_reg(110) <= "00010101000101100000000100100001";
                        f_reg(111) <= "10101100000010000000010001001000";
                        f_reg(112) <= "00000001000000010110000000000100";
                        f_reg(113) <= "00000010110011111101000000000100";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00000000000000000000000000000000";
                        f_reg(116) <= "00000001100010110110100000101011";
                        f_reg(117) <= "00000011010110011101100000101011";
                        f_reg(118) <= "00000000000010000111000110000010";
                        f_reg(119) <= "00000000000101101110000110000010";
                        f_reg(120) <= "00010100001011110000000100010111";
                        f_reg(121) <= "10101100000000010000010001001100";
                        f_reg(122) <= "00000001001001010010100000101011";
                        f_reg(123) <= "00000010111100111001100000101011";
                        f_reg(124) <= "00000000001001100001000000100011";
                        f_reg(125) <= "00000001111101001000000000100011";
                        f_reg(126) <= "00000000100000110011100000100100";
                        f_reg(127) <= "00000010010100011010100000100100";
                        f_reg(128) <= "00101001110000111000100100101101";
                        f_reg(129) <= "00101011100100011000100100101101";
                        f_reg(130) <= "00010100011100010000000100001101";
                        f_reg(131) <= "10101100000000110000010001111100";
                        f_reg(132) <= "00000000100001100001100000100111";
                        f_reg(133) <= "00000010010101001000100000100111";
                        f_reg(134) <= "00010100011100010000000100001001";
                        f_reg(135) <= "10101100000000110000010010000000";
                        f_reg(136) <= "00101101000000110100100000000010";
                        f_reg(137) <= "00101110110100010100100000000010";
                        f_reg(138) <= "00010100011100010000000100000101";
                        f_reg(139) <= "10101100000000110000010010000100";
                        f_reg(140) <= "00000001101000010001100000100100";
                        f_reg(141) <= "00000011011011111000100000100100";
                        f_reg(142) <= "00010101100110100000000100000001";
                        f_reg(143) <= "10101100000011000000010001010000";
                        f_reg(144) <= "00000000000000010110000000000110";
                        f_reg(145) <= "00000000000011111101000000000110";
                        f_reg(146) <= "10001100000000010000010010000000";
                        f_reg(147) <= "10001100000011110000010010000000";
                        f_reg(148) <= "00010100001011111111111111111110";
                        f_reg(149) <= "00010101000101100000000011111010";
                        f_reg(150) <= "10101100000010000000010010000000";
                        f_reg(151) <= "00000000001011100100000000100001";
                        f_reg(152) <= "00000001111111001011000000100001";
                        f_reg(153) <= "00000000101000100111000000101010";
                        f_reg(154) <= "00000010011100001110000000101010";
                        f_reg(155) <= "00000001011010100001000000100001";
                        f_reg(156) <= "00000011001110001000000000100001";
                        f_reg(157) <= "00010101010110000000000011110010";
                        f_reg(158) <= "10101100000010100000010001010100";
                        f_reg(159) <= "00000000000000000000000000000000";
                        f_reg(160) <= "00000000000000000000000000000000";
                        f_reg(161) <= "10001100000010100000010010000100";
                        f_reg(162) <= "10001100000110000000010010000100";
                        f_reg(163) <= "00010101010110001111111111111110";
                        f_reg(164) <= "00010101000101100000000011101011";
                        f_reg(165) <= "10101100000010000000010010000100";
                        f_reg(166) <= "00000001010000010100000000100101";
                        f_reg(167) <= "00000011000011111011000000100101";
                        f_reg(168) <= "00010101010110000000000011100111";
                        f_reg(169) <= "10101100000010100000010010001000";
                        f_reg(170) <= "00000000000010010101010000000011";
                        f_reg(171) <= "00000000000101111100010000000011";
                        f_reg(172) <= "00010101000101100000000011100011";
                        f_reg(173) <= "10101100000010000000010001011000";
                        f_reg(174) <= "00000000110001000011000000100010";
                        f_reg(175) <= "00000010100100101010000000100010";
                        f_reg(176) <= "00100101110010011101010011110111";
                        f_reg(177) <= "00100111100101111101010011110111";
                        f_reg(178) <= "00000000101011010010100000100111";
                        f_reg(179) <= "00000010011110111001100000100111";
                        f_reg(180) <= "00000000000010000010010000000011";
                        f_reg(181) <= "00000000000101101001010000000011";
                        f_reg(182) <= "00101101011011100001011001001101";
                        f_reg(183) <= "00101111001111000001011001001101";
                        f_reg(184) <= "00000001001001110110100000101011";
                        f_reg(185) <= "00000010111101011101100000101011";
                        f_reg(186) <= "00000000010000010101100000100000";
                        f_reg(187) <= "00000010000011111100100000100000";
                        f_reg(188) <= "00000000011000000100100000100100";
                        f_reg(189) <= "00000010001000001011100000100100";
                        f_reg(190) <= "00010101001101110000000011010001";
                        f_reg(191) <= "10101100000010010000010001011100";
                        f_reg(192) <= "00110001100001111000000001111000";
                        f_reg(193) <= "00110011010101011000000001111000";
                        f_reg(194) <= "00000001011011010001000000100011";
                        f_reg(195) <= "00000011001110111000000000100011";
                        f_reg(196) <= "00000001010001000000100000100010";
                        f_reg(197) <= "00000011000100100111100000100010";
                        f_reg(198) <= "00000000110011010001100000101011";
                        f_reg(199) <= "00000010100110111000100000101011";
                        f_reg(200) <= "10001100000010010000010010000000";
                        f_reg(201) <= "10001100000101110000010010000000";
                        f_reg(202) <= "00010101001101111111111111111110";
                        f_reg(203) <= "00000001011010010110000000100101";
                        f_reg(204) <= "00000011001101111101000000100101";
                        f_reg(205) <= "00100101000010101000000100111100";
                        f_reg(206) <= "00100110110110001000000100111100";
                        f_reg(207) <= "00111000101001001100000101001101";
                        f_reg(208) <= "00111010011100101100000101001101";
                        f_reg(209) <= "10001100000010110000010001111100";
                        f_reg(210) <= "10001100000110010000010001111100";
                        f_reg(211) <= "00010101011110011111111111111110";
                        f_reg(212) <= "00010101011110010000000010111011";
                        f_reg(213) <= "10101100000010110000010001100000";
                        f_reg(214) <= "00101100011010010110110111011111";
                        f_reg(215) <= "00101110001101110110110111011111";
                        f_reg(216) <= "00010101100110100000000010110111";
                        f_reg(217) <= "10101100000011000000010001100100";
                        f_reg(218) <= "00010101010110000000000010110101";
                        f_reg(219) <= "10101100000010100000010001101000";
                        f_reg(220) <= "00000001101001000100000000000100";
                        f_reg(221) <= "00000011011100101011000000000100";
                        f_reg(222) <= "00000000111011100010100000101010";
                        f_reg(223) <= "00000010101111001001100000101010";
                        f_reg(224) <= "00000000001010010101100000100110";
                        f_reg(225) <= "00000001111101111100100000100110";
                        f_reg(226) <= "00000000110000110110000000100111";
                        f_reg(227) <= "00000010100100011101000000100111";
                        f_reg(228) <= "00000000000000000000000000000000";
                        f_reg(229) <= "00000000000000000000000000000000";
                        f_reg(230) <= "00010101100110100000000010101001";
                        f_reg(231) <= "10101100000011000000010001101100";
                        f_reg(232) <= "00010100101100110000000010100111";
                        f_reg(233) <= "10101100000001010000010001110000";
                        f_reg(234) <= "00000001000000000101000000100100";
                        f_reg(235) <= "00000010110000001100000000100100";
                        f_reg(236) <= "10001100000001000000010010001000";
                        f_reg(237) <= "10001100000100100000010010001000";
                        f_reg(238) <= "00010100100100101111111111111110";
                        f_reg(239) <= "00000000100000100110100000100010";
                        f_reg(240) <= "00000010010100001101100000100010";
                        f_reg(241) <= "10001100000001110000010010000100";
                        f_reg(242) <= "10001100000101010000010010000100";
                        f_reg(243) <= "00010100111101011111111111111110";
                        f_reg(244) <= "00000000111010110111000000100000";
                        f_reg(245) <= "00000010101110011110000000100000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00110101010000010111000001000101";
                        f_reg(249) <= "00110111000011110111000001000101";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00000000000000000000000000000000";
                        f_reg(252) <= "00000000001011010100100000101011";
                        f_reg(253) <= "00000001111110111011100000101011";
                        f_reg(254) <= "00010101001101110000000010010001";
                        f_reg(255) <= "10101100000010010000010001110100";
                        f_reg(256) <= "00000000000011100111001111000000";
                        f_reg(257) <= "00000000000111001110001111000000";
                        f_reg(258) <= "00000000000000000000000000000000";
                        f_reg(259) <= "00000000000000000000000000000000";
                        f_reg(260) <= "00010101110111000000000010001011";
                        f_reg(261) <= "10101100000011100000010001111000";
                        f_reg(262) <= "00100011110111011111111100000110";
                        f_reg(263) <= "00010011101000000000000000011101";
                        f_reg(264) <= "00100011110111011111111000001100";
                        f_reg(265) <= "00010011101000000000000000011011";
                        f_reg(266) <= "00100011110111011111110100010010";
                        f_reg(267) <= "00010011101000000000000000011001";
                        f_reg(268) <= "00100011110111101111111111111111";
                        f_reg(269) <= "00100011111111111111111111111111";
                        f_reg(270) <= "00010111110111110000000010000001";
                        f_reg(271) <= "00011111111000001111111101000101";
                        f_reg(272) <= "00010000000000000000000100001100";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "00000000000000000000000000000000";
                        f_reg(287) <= "00000000000000000000000000000000";
                        f_reg(288) <= "00000000000000000000000000000000";
                        f_reg(289) <= "00000000000000000000000000000000";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "10001100000111010000011111100000";
                        f_reg(293) <= "00011111101000000000000000000011";
                        f_reg(294) <= "00100000000111010000000000111100";
                        f_reg(295) <= "00010000000000000000000000000010";
                        f_reg(296) <= "00100000000111010000000000000000";
                        f_reg(297) <= "00010100001011110000000001100110";
                        f_reg(298) <= "10101111101000010000011101101000";
                        f_reg(299) <= "10001100000111010000011111100000";
                        f_reg(300) <= "00011111101000000000000000000011";
                        f_reg(301) <= "00100000000111010000000000111100";
                        f_reg(302) <= "00010000000000000000000000000010";
                        f_reg(303) <= "00100000000111010000000000000000";
                        f_reg(304) <= "00010100010100000000000001011111";
                        f_reg(305) <= "10101111101000100000011101101100";
                        f_reg(306) <= "10001100000111010000011111100000";
                        f_reg(307) <= "00011111101000000000000000000011";
                        f_reg(308) <= "00100000000111010000000000111100";
                        f_reg(309) <= "00010000000000000000000000000010";
                        f_reg(310) <= "00100000000111010000000000000000";
                        f_reg(311) <= "00010100011100010000000001011000";
                        f_reg(312) <= "10101111101000110000011101110000";
                        f_reg(313) <= "10001100000111010000011111100000";
                        f_reg(314) <= "00011111101000000000000000000011";
                        f_reg(315) <= "00100000000111010000000000111100";
                        f_reg(316) <= "00010000000000000000000000000010";
                        f_reg(317) <= "00100000000111010000000000000000";
                        f_reg(318) <= "00010100100100100000000001010001";
                        f_reg(319) <= "10101111101001000000011101110100";
                        f_reg(320) <= "10001100000111010000011111100000";
                        f_reg(321) <= "00011111101000000000000000000011";
                        f_reg(322) <= "00100000000111010000000000111100";
                        f_reg(323) <= "00010000000000000000000000000010";
                        f_reg(324) <= "00100000000111010000000000000000";
                        f_reg(325) <= "00010100101100110000000001001010";
                        f_reg(326) <= "10101111101001010000011101111000";
                        f_reg(327) <= "10001100000111010000011111100000";
                        f_reg(328) <= "00011111101000000000000000000011";
                        f_reg(329) <= "00100000000111010000000000111100";
                        f_reg(330) <= "00010000000000000000000000000010";
                        f_reg(331) <= "00100000000111010000000000000000";
                        f_reg(332) <= "00010100110101000000000001000011";
                        f_reg(333) <= "10101111101001100000011101111100";
                        f_reg(334) <= "10001100000111010000011111100000";
                        f_reg(335) <= "00011111101000000000000000000011";
                        f_reg(336) <= "00100000000111010000000000111100";
                        f_reg(337) <= "00010000000000000000000000000010";
                        f_reg(338) <= "00100000000111010000000000000000";
                        f_reg(339) <= "00010100111101010000000000111100";
                        f_reg(340) <= "10101111101001110000011110000000";
                        f_reg(341) <= "10001100000111010000011111100000";
                        f_reg(342) <= "00011111101000000000000000000011";
                        f_reg(343) <= "00100000000111010000000000111100";
                        f_reg(344) <= "00010000000000000000000000000010";
                        f_reg(345) <= "00100000000111010000000000000000";
                        f_reg(346) <= "00010101000101100000000000110101";
                        f_reg(347) <= "10101111101010000000011110000100";
                        f_reg(348) <= "10001100000111010000011111100000";
                        f_reg(349) <= "00011111101000000000000000000011";
                        f_reg(350) <= "00100000000111010000000000111100";
                        f_reg(351) <= "00010000000000000000000000000010";
                        f_reg(352) <= "00100000000111010000000000000000";
                        f_reg(353) <= "00010101001101110000000000101110";
                        f_reg(354) <= "10101111101010010000011110001000";
                        f_reg(355) <= "10001100000111010000011111100000";
                        f_reg(356) <= "00011111101000000000000000000011";
                        f_reg(357) <= "00100000000111010000000000111100";
                        f_reg(358) <= "00010000000000000000000000000010";
                        f_reg(359) <= "00100000000111010000000000000000";
                        f_reg(360) <= "00010101010110000000000000100111";
                        f_reg(361) <= "10101111101010100000011110001100";
                        f_reg(362) <= "10001100000111010000011111100000";
                        f_reg(363) <= "00011111101000000000000000000011";
                        f_reg(364) <= "00100000000111010000000000111100";
                        f_reg(365) <= "00010000000000000000000000000010";
                        f_reg(366) <= "00100000000111010000000000000000";
                        f_reg(367) <= "00010101011110010000000000100000";
                        f_reg(368) <= "10101111101010110000011110010000";
                        f_reg(369) <= "10001100000111010000011111100000";
                        f_reg(370) <= "00011111101000000000000000000011";
                        f_reg(371) <= "00100000000111010000000000111100";
                        f_reg(372) <= "00010000000000000000000000000010";
                        f_reg(373) <= "00100000000111010000000000000000";
                        f_reg(374) <= "00010101100110100000000000011001";
                        f_reg(375) <= "10101111101011000000011110010100";
                        f_reg(376) <= "10001100000111010000011111100000";
                        f_reg(377) <= "00011111101000000000000000000011";
                        f_reg(378) <= "00100000000111010000000000111100";
                        f_reg(379) <= "00010000000000000000000000000010";
                        f_reg(380) <= "00100000000111010000000000000000";
                        f_reg(381) <= "00010101101110110000000000010010";
                        f_reg(382) <= "10101111101011010000011110011000";
                        f_reg(383) <= "10001100000111010000011111100000";
                        f_reg(384) <= "00011111101000000000000000000011";
                        f_reg(385) <= "00100000000111010000000000111100";
                        f_reg(386) <= "00010000000000000000000000000010";
                        f_reg(387) <= "00100000000111010000000000000000";
                        f_reg(388) <= "00010101110111000000000000001011";
                        f_reg(389) <= "10101111101011100000011110011100";
                        f_reg(390) <= "10001100000111010000011111100000";
                        f_reg(391) <= "00011111101000000000000000000011";
                        f_reg(392) <= "00100000000111010000000000111100";
                        f_reg(393) <= "00010000000000000000000000000010";
                        f_reg(394) <= "00100000000111010000000000000000";
                        f_reg(395) <= "00010111110111110000000000000100";
                        f_reg(396) <= "10101111101111100000011110100000";
                        f_reg(397) <= "10101100000111010000011111100000";
                        f_reg(398) <= "00010000000000001111111101111110";
                        f_reg(399) <= "10001100000111010000011111100000";
                        f_reg(400) <= "10001111101000010000011101101000";
                        f_reg(401) <= "10001100000111010000011111100000";
                        f_reg(402) <= "10001111101011110000011101101000";
                        f_reg(403) <= "00010100001011111111111111111100";
                        f_reg(404) <= "10001100000111010000011111100000";
                        f_reg(405) <= "10001111101000100000011101101100";
                        f_reg(406) <= "10001100000111010000011111100000";
                        f_reg(407) <= "10001111101100000000011101101100";
                        f_reg(408) <= "00010100010100001111111111111100";
                        f_reg(409) <= "10001100000111010000011111100000";
                        f_reg(410) <= "10001111101000110000011101110000";
                        f_reg(411) <= "10001100000111010000011111100000";
                        f_reg(412) <= "10001111101100010000011101110000";
                        f_reg(413) <= "00010100011100011111111111111100";
                        f_reg(414) <= "10001100000111010000011111100000";
                        f_reg(415) <= "10001111101001000000011101110100";
                        f_reg(416) <= "10001100000111010000011111100000";
                        f_reg(417) <= "10001111101100100000011101110100";
                        f_reg(418) <= "00010100100100101111111111111100";
                        f_reg(419) <= "10001100000111010000011111100000";
                        f_reg(420) <= "10001111101001010000011101111000";
                        f_reg(421) <= "10001100000111010000011111100000";
                        f_reg(422) <= "10001111101100110000011101111000";
                        f_reg(423) <= "00010100101100111111111111111100";
                        f_reg(424) <= "10001100000111010000011111100000";
                        f_reg(425) <= "10001111101001100000011101111100";
                        f_reg(426) <= "10001100000111010000011111100000";
                        f_reg(427) <= "10001111101101000000011101111100";
                        f_reg(428) <= "00010100110101001111111111111100";
                        f_reg(429) <= "10001100000111010000011111100000";
                        f_reg(430) <= "10001111101001110000011110000000";
                        f_reg(431) <= "10001100000111010000011111100000";
                        f_reg(432) <= "10001111101101010000011110000000";
                        f_reg(433) <= "00010100111101011111111111111100";
                        f_reg(434) <= "10001100000111010000011111100000";
                        f_reg(435) <= "10001111101010000000011110000100";
                        f_reg(436) <= "10001100000111010000011111100000";
                        f_reg(437) <= "10001111101101100000011110000100";
                        f_reg(438) <= "00010101000101101111111111111100";
                        f_reg(439) <= "10001100000111010000011111100000";
                        f_reg(440) <= "10001111101010010000011110001000";
                        f_reg(441) <= "10001100000111010000011111100000";
                        f_reg(442) <= "10001111101101110000011110001000";
                        f_reg(443) <= "00010101001101111111111111111100";
                        f_reg(444) <= "10001100000111010000011111100000";
                        f_reg(445) <= "10001111101010100000011110001100";
                        f_reg(446) <= "10001100000111010000011111100000";
                        f_reg(447) <= "10001111101110000000011110001100";
                        f_reg(448) <= "00010101010110001111111111111100";
                        f_reg(449) <= "10001100000111010000011111100000";
                        f_reg(450) <= "10001111101010110000011110010000";
                        f_reg(451) <= "10001100000111010000011111100000";
                        f_reg(452) <= "10001111101110010000011110010000";
                        f_reg(453) <= "00010101011110011111111111111100";
                        f_reg(454) <= "10001100000111010000011111100000";
                        f_reg(455) <= "10001111101011000000011110010100";
                        f_reg(456) <= "10001100000111010000011111100000";
                        f_reg(457) <= "10001111101110100000011110010100";
                        f_reg(458) <= "00010101100110101111111111111100";
                        f_reg(459) <= "10001100000111010000011111100000";
                        f_reg(460) <= "10001111101011010000011110011000";
                        f_reg(461) <= "10001100000111010000011111100000";
                        f_reg(462) <= "10001111101110110000011110011000";
                        f_reg(463) <= "00010101101110111111111111111100";
                        f_reg(464) <= "10001100000111010000011111100000";
                        f_reg(465) <= "10001111101011100000011110011100";
                        f_reg(466) <= "10001100000111010000011111100000";
                        f_reg(467) <= "10001111101111000000011110011100";
                        f_reg(468) <= "00010101110111001111111111111100";
                        f_reg(469) <= "10001100000111010000011111100000";
                        f_reg(470) <= "10001111101111100000011110100000";
                        f_reg(471) <= "10001100000111010000011111100000";
                        f_reg(472) <= "10001111101111110000011110100000";
                        f_reg(473) <= "00010111110111111111111111111100";
                        f_reg(474) <= "00010000000000001111111100110010";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000001111100111";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010001001011010101";
                        f_reg(4) <= "00000000001000010001000000100010";
                        f_reg(5) <= "00101000001000110010100010011111";
                        f_reg(6) <= "00000000001000010010000000100000";
                        f_reg(7) <= "00000000000000100010100001000011";
                        f_reg(8) <= "00000000101000110011000000100011";
                        f_reg(9) <= "00000000010000100011100000100101";
                        f_reg(10) <= "00000000000000000100000111000011";
                        f_reg(11) <= "10101100000010000000010001000000";
                        f_reg(12) <= "10101100000000010000010001000100";
                        f_reg(13) <= "00000000100001000100100000000110";
                        f_reg(14) <= "00000000111001110101000000101011";
                        f_reg(15) <= "00000000110010100101100000100111";
                        f_reg(16) <= "10101100000010000000010001001000";
                        f_reg(17) <= "00000001000000010110000000000100";
                        f_reg(18) <= "00000000000000000000000000000000";
                        f_reg(19) <= "00000001100010110110100000101011";
                        f_reg(20) <= "00000000000010000111000110000010";
                        f_reg(21) <= "10101100000000010000010001001100";
                        f_reg(22) <= "00000001001001010010100000101011";
                        f_reg(23) <= "00000000001001100111100000100011";
                        f_reg(24) <= "00000000100000111000000000100100";
                        f_reg(25) <= "00101001110100011000100100101101";
                        f_reg(26) <= "00000000100001101001000000100111";
                        f_reg(27) <= "00101101000100110100100000000010";
                        f_reg(28) <= "00000001101000011010000000100100";
                        f_reg(29) <= "10101100000011000000010001010000";
                        f_reg(30) <= "00000000000000011010100000000110";
                        f_reg(31) <= "00000010010011101011000000100001";
                        f_reg(32) <= "00000000101011111011100000101010";
                        f_reg(33) <= "00000001011010101100000000100001";
                        f_reg(34) <= "10101100000010100000010001010100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000010011100101100100000100101";
                        f_reg(37) <= "00000000000010011101010000000011";
                        f_reg(38) <= "10101100000110010000010001011000";
                        f_reg(39) <= "00000000110001000011000000100010";
                        f_reg(40) <= "00100110111110111101010011110111";
                        f_reg(41) <= "00000000101011010010100000100111";
                        f_reg(42) <= "00000000000110011110010000000011";
                        f_reg(43) <= "00101101011111010001011001001101";
                        f_reg(44) <= "00000011011100001111000000101011";
                        f_reg(45) <= "00000011000100100001000000100000";
                        f_reg(46) <= "00000010100000000011100000100100";
                        f_reg(47) <= "10101100000001110000010001011100";
                        f_reg(48) <= "00110010101000111000000001111000";
                        f_reg(49) <= "00000000010111100110000000100011";
                        f_reg(50) <= "00000011010111000000100000100010";
                        f_reg(51) <= "00000000110111100111000000101011";
                        f_reg(52) <= "00000000010010000111100000100101";
                        f_reg(53) <= "00100111001010101000000100111100";
                        f_reg(54) <= "00111000101010011100000101001101";
                        f_reg(55) <= "10101100000100010000010001100000";
                        f_reg(56) <= "00101101110001000110110111011111";
                        f_reg(57) <= "10101100000011110000010001100100";
                        f_reg(58) <= "10101100000010100000010001101000";
                        f_reg(59) <= "00000011110010011011100000000100";
                        f_reg(60) <= "00000000011111010110100000101010";
                        f_reg(61) <= "00000000001001000101100000100110";
                        f_reg(62) <= "00000000110011101101100000100111";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000110110000010001101100";
                        f_reg(65) <= "10101100000011010000010001110000";
                        f_reg(66) <= "00000010111000001000000000100100";
                        f_reg(67) <= "00000010011011001100000000100010";
                        f_reg(68) <= "00000010110010111001000000100000";
                        f_reg(69) <= "00000000000000000000000000000000";
                        f_reg(70) <= "00110110000101000111000001000101";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000010100110000011100000101011";
                        f_reg(73) <= "10101100000001110000010001110100";
                        f_reg(74) <= "00000000000100101001001111000000";
                        f_reg(75) <= "00000000000000000000000000000000";
                        f_reg(76) <= "10101100000100100000010001111000";
                        f_reg(77) <= "00100011111111111111111111111111";
                        f_reg(78) <= "00011111111000001111111110110101";
                        f_reg(79) <= "00010000000000000000000111001101";
                        f_reg(80) <= "00111100000111100000001111100111";
                        f_reg(81) <= "00111100000111110000001111100111";
                        f_reg(82) <= "00000000000111101111010000000010";
                        f_reg(83) <= "00000000000111111111110000000010";
                        f_reg(84) <= "00111100000000010001001011010101";
                        f_reg(85) <= "00111100000011110001001011010101";
                        f_reg(86) <= "00000000001000010001000000100010";
                        f_reg(87) <= "00000001111011111000000000100010";
                        f_reg(88) <= "00101000001000110010100010011111";
                        f_reg(89) <= "00101001111100010010100010011111";
                        f_reg(90) <= "00000000001000010010000000100000";
                        f_reg(91) <= "00000001111011111001000000100000";
                        f_reg(92) <= "00000000000000100010100001000011";
                        f_reg(93) <= "00000000000100001001100001000011";
                        f_reg(94) <= "00000000101000110011000000100011";
                        f_reg(95) <= "00000010011100011010000000100011";
                        f_reg(96) <= "00000000010000100011100000100101";
                        f_reg(97) <= "00000010000100001010100000100101";
                        f_reg(98) <= "00000000000000000100000111000011";
                        f_reg(99) <= "00000000000000001011000111000011";
                        f_reg(100) <= "00010101000101100000000100101011";
                        f_reg(101) <= "10101100000010000000010001000000";
                        f_reg(102) <= "00010100001011110000000100101001";
                        f_reg(103) <= "10101100000000010000010001000100";
                        f_reg(104) <= "00000000100001000100100000000110";
                        f_reg(105) <= "00000010010100101011100000000110";
                        f_reg(106) <= "00000000111001110101000000101011";
                        f_reg(107) <= "00000010101101011100000000101011";
                        f_reg(108) <= "00000000110010100101100000100111";
                        f_reg(109) <= "00000010100110001100100000100111";
                        f_reg(110) <= "00010101000101100000000100100001";
                        f_reg(111) <= "10101100000010000000010001001000";
                        f_reg(112) <= "00000001000000010110000000000100";
                        f_reg(113) <= "00000010110011111101000000000100";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00000000000000000000000000000000";
                        f_reg(116) <= "00000001100010110110100000101011";
                        f_reg(117) <= "00000011010110011101100000101011";
                        f_reg(118) <= "00000000000010000111000110000010";
                        f_reg(119) <= "00000000000101101110000110000010";
                        f_reg(120) <= "00010100001011110000000100010111";
                        f_reg(121) <= "10101100000000010000010001001100";
                        f_reg(122) <= "00000001001001010010100000101011";
                        f_reg(123) <= "00000010111100111001100000101011";
                        f_reg(124) <= "00000000001001100001000000100011";
                        f_reg(125) <= "00000001111101001000000000100011";
                        f_reg(126) <= "00000000100000110011100000100100";
                        f_reg(127) <= "00000010010100011010100000100100";
                        f_reg(128) <= "00101001110000111000100100101101";
                        f_reg(129) <= "00101011100100011000100100101101";
                        f_reg(130) <= "00010100011100010000000100001101";
                        f_reg(131) <= "10101100000000110000010001111100";
                        f_reg(132) <= "00000000100001100001100000100111";
                        f_reg(133) <= "00000010010101001000100000100111";
                        f_reg(134) <= "00010100011100010000000100001001";
                        f_reg(135) <= "10101100000000110000010010000000";
                        f_reg(136) <= "00101101000000110100100000000010";
                        f_reg(137) <= "00101110110100010100100000000010";
                        f_reg(138) <= "00010100011100010000000100000101";
                        f_reg(139) <= "10101100000000110000010010000100";
                        f_reg(140) <= "00000001101000010001100000100100";
                        f_reg(141) <= "00000011011011111000100000100100";
                        f_reg(142) <= "00010101100110100000000100000001";
                        f_reg(143) <= "10101100000011000000010001010000";
                        f_reg(144) <= "00000000000000010110000000000110";
                        f_reg(145) <= "00000000000011111101000000000110";
                        f_reg(146) <= "10001100000000010000010010000000";
                        f_reg(147) <= "10001100000011110000010010000000";
                        f_reg(148) <= "00010100001011111111111111111110";
                        f_reg(149) <= "00010101000101100000000011111010";
                        f_reg(150) <= "10101100000010000000010010000000";
                        f_reg(151) <= "00000000001011100100000000100001";
                        f_reg(152) <= "00000001111111001011000000100001";
                        f_reg(153) <= "00000000101000100111000000101010";
                        f_reg(154) <= "00000010011100001110000000101010";
                        f_reg(155) <= "00000001011010100001000000100001";
                        f_reg(156) <= "00000011001110001000000000100001";
                        f_reg(157) <= "00010101010110000000000011110010";
                        f_reg(158) <= "10101100000010100000010001010100";
                        f_reg(159) <= "00000000000000000000000000000000";
                        f_reg(160) <= "00000000000000000000000000000000";
                        f_reg(161) <= "10001100000010100000010010000100";
                        f_reg(162) <= "10001100000110000000010010000100";
                        f_reg(163) <= "00010101010110001111111111111110";
                        f_reg(164) <= "00010101000101100000000011101011";
                        f_reg(165) <= "10101100000010000000010010000100";
                        f_reg(166) <= "00000001010000010100000000100101";
                        f_reg(167) <= "00000011000011111011000000100101";
                        f_reg(168) <= "00010101010110000000000011100111";
                        f_reg(169) <= "10101100000010100000010010001000";
                        f_reg(170) <= "00000000000010010101010000000011";
                        f_reg(171) <= "00000000000101111100010000000011";
                        f_reg(172) <= "00010101000101100000000011100011";
                        f_reg(173) <= "10101100000010000000010001011000";
                        f_reg(174) <= "00000000110001000011000000100010";
                        f_reg(175) <= "00000010100100101010000000100010";
                        f_reg(176) <= "00100101110010011101010011110111";
                        f_reg(177) <= "00100111100101111101010011110111";
                        f_reg(178) <= "00000000101011010010100000100111";
                        f_reg(179) <= "00000010011110111001100000100111";
                        f_reg(180) <= "00000000000010000010010000000011";
                        f_reg(181) <= "00000000000101101001010000000011";
                        f_reg(182) <= "00101101011011100001011001001101";
                        f_reg(183) <= "00101111001111000001011001001101";
                        f_reg(184) <= "00000001001001110110100000101011";
                        f_reg(185) <= "00000010111101011101100000101011";
                        f_reg(186) <= "00000000010000010101100000100000";
                        f_reg(187) <= "00000010000011111100100000100000";
                        f_reg(188) <= "00000000011000000100100000100100";
                        f_reg(189) <= "00000010001000001011100000100100";
                        f_reg(190) <= "00010101001101110000000011010001";
                        f_reg(191) <= "10101100000010010000010001011100";
                        f_reg(192) <= "00110001100001111000000001111000";
                        f_reg(193) <= "00110011010101011000000001111000";
                        f_reg(194) <= "00000001011011010001000000100011";
                        f_reg(195) <= "00000011001110111000000000100011";
                        f_reg(196) <= "00000001010001000000100000100010";
                        f_reg(197) <= "00000011000100100111100000100010";
                        f_reg(198) <= "00000000110011010001100000101011";
                        f_reg(199) <= "00000010100110111000100000101011";
                        f_reg(200) <= "10001100000010010000010010000000";
                        f_reg(201) <= "10001100000101110000010010000000";
                        f_reg(202) <= "00010101001101111111111111111110";
                        f_reg(203) <= "00000001011010010110000000100101";
                        f_reg(204) <= "00000011001101111101000000100101";
                        f_reg(205) <= "00100101000010101000000100111100";
                        f_reg(206) <= "00100110110110001000000100111100";
                        f_reg(207) <= "00111000101001001100000101001101";
                        f_reg(208) <= "00111010011100101100000101001101";
                        f_reg(209) <= "10001100000010110000010001111100";
                        f_reg(210) <= "10001100000110010000010001111100";
                        f_reg(211) <= "00010101011110011111111111111110";
                        f_reg(212) <= "00010101011110010000000010111011";
                        f_reg(213) <= "10101100000010110000010001100000";
                        f_reg(214) <= "00101100011010010110110111011111";
                        f_reg(215) <= "00101110001101110110110111011111";
                        f_reg(216) <= "00010101100110100000000010110111";
                        f_reg(217) <= "10101100000011000000010001100100";
                        f_reg(218) <= "00010101010110000000000010110101";
                        f_reg(219) <= "10101100000010100000010001101000";
                        f_reg(220) <= "00000001101001000100000000000100";
                        f_reg(221) <= "00000011011100101011000000000100";
                        f_reg(222) <= "00000000111011100010100000101010";
                        f_reg(223) <= "00000010101111001001100000101010";
                        f_reg(224) <= "00000000001010010101100000100110";
                        f_reg(225) <= "00000001111101111100100000100110";
                        f_reg(226) <= "00000000110000110110000000100111";
                        f_reg(227) <= "00000010100100011101000000100111";
                        f_reg(228) <= "00000000000000000000000000000000";
                        f_reg(229) <= "00000000000000000000000000000000";
                        f_reg(230) <= "00010101100110100000000010101001";
                        f_reg(231) <= "10101100000011000000010001101100";
                        f_reg(232) <= "00010100101100110000000010100111";
                        f_reg(233) <= "10101100000001010000010001110000";
                        f_reg(234) <= "00000001000000000101000000100100";
                        f_reg(235) <= "00000010110000001100000000100100";
                        f_reg(236) <= "10001100000001000000010010001000";
                        f_reg(237) <= "10001100000100100000010010001000";
                        f_reg(238) <= "00010100100100101111111111111110";
                        f_reg(239) <= "00000000100000100110100000100010";
                        f_reg(240) <= "00000010010100001101100000100010";
                        f_reg(241) <= "10001100000001110000010010000100";
                        f_reg(242) <= "10001100000101010000010010000100";
                        f_reg(243) <= "00010100111101011111111111111110";
                        f_reg(244) <= "00000000111010110111000000100000";
                        f_reg(245) <= "00000010101110011110000000100000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00110101010000010111000001000101";
                        f_reg(249) <= "00110111000011110111000001000101";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00000000000000000000000000000000";
                        f_reg(252) <= "00000000001011010100100000101011";
                        f_reg(253) <= "00000001111110111011100000101011";
                        f_reg(254) <= "00010101001101110000000010010001";
                        f_reg(255) <= "10101100000010010000010001110100";
                        f_reg(256) <= "00000000000011100111001111000000";
                        f_reg(257) <= "00000000000111001110001111000000";
                        f_reg(258) <= "00000000000000000000000000000000";
                        f_reg(259) <= "00000000000000000000000000000000";
                        f_reg(260) <= "00010101110111000000000010001011";
                        f_reg(261) <= "10101100000011100000010001111000";
                        f_reg(262) <= "00100011110111011111111100000110";
                        f_reg(263) <= "00010011101000000000000000011101";
                        f_reg(264) <= "00100011110111011111111000001100";
                        f_reg(265) <= "00010011101000000000000000011011";
                        f_reg(266) <= "00100011110111011111110100010010";
                        f_reg(267) <= "00010011101000000000000000011001";
                        f_reg(268) <= "00100011110111101111111111111111";
                        f_reg(269) <= "00100011111111111111111111111111";
                        f_reg(270) <= "00010111110111110000000010000001";
                        f_reg(271) <= "00011111111000001111111101000101";
                        f_reg(272) <= "00010000000000000000000100001100";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "00000000000000000000000000000000";
                        f_reg(287) <= "00000000000000000000000000000000";
                        f_reg(288) <= "00000000000000000000000000000000";
                        f_reg(289) <= "00000000000000000000000000000000";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "10001100000111010000011111100000";
                        f_reg(293) <= "00011111101000000000000000000011";
                        f_reg(294) <= "00100000000111010000000000111100";
                        f_reg(295) <= "00010000000000000000000000000010";
                        f_reg(296) <= "00100000000111010000000000000000";
                        f_reg(297) <= "00010100001011110000000001100110";
                        f_reg(298) <= "10101111101000010000011101101000";
                        f_reg(299) <= "10001100000111010000011111100000";
                        f_reg(300) <= "00011111101000000000000000000011";
                        f_reg(301) <= "00100000000111010000000000111100";
                        f_reg(302) <= "00010000000000000000000000000010";
                        f_reg(303) <= "00100000000111010000000000000000";
                        f_reg(304) <= "00010100010100000000000001011111";
                        f_reg(305) <= "10101111101000100000011101101100";
                        f_reg(306) <= "10001100000111010000011111100000";
                        f_reg(307) <= "00011111101000000000000000000011";
                        f_reg(308) <= "00100000000111010000000000111100";
                        f_reg(309) <= "00010000000000000000000000000010";
                        f_reg(310) <= "00100000000111010000000000000000";
                        f_reg(311) <= "00010100011100010000000001011000";
                        f_reg(312) <= "10101111101000110000011101110000";
                        f_reg(313) <= "10001100000111010000011111100000";
                        f_reg(314) <= "00011111101000000000000000000011";
                        f_reg(315) <= "00100000000111010000000000111100";
                        f_reg(316) <= "00010000000000000000000000000010";
                        f_reg(317) <= "00100000000111010000000000000000";
                        f_reg(318) <= "00010100100100100000000001010001";
                        f_reg(319) <= "10101111101001000000011101110100";
                        f_reg(320) <= "10001100000111010000011111100000";
                        f_reg(321) <= "00011111101000000000000000000011";
                        f_reg(322) <= "00100000000111010000000000111100";
                        f_reg(323) <= "00010000000000000000000000000010";
                        f_reg(324) <= "00100000000111010000000000000000";
                        f_reg(325) <= "00010100101100110000000001001010";
                        f_reg(326) <= "10101111101001010000011101111000";
                        f_reg(327) <= "10001100000111010000011111100000";
                        f_reg(328) <= "00011111101000000000000000000011";
                        f_reg(329) <= "00100000000111010000000000111100";
                        f_reg(330) <= "00010000000000000000000000000010";
                        f_reg(331) <= "00100000000111010000000000000000";
                        f_reg(332) <= "00010100110101000000000001000011";
                        f_reg(333) <= "10101111101001100000011101111100";
                        f_reg(334) <= "10001100000111010000011111100000";
                        f_reg(335) <= "00011111101000000000000000000011";
                        f_reg(336) <= "00100000000111010000000000111100";
                        f_reg(337) <= "00010000000000000000000000000010";
                        f_reg(338) <= "00100000000111010000000000000000";
                        f_reg(339) <= "00010100111101010000000000111100";
                        f_reg(340) <= "10101111101001110000011110000000";
                        f_reg(341) <= "10001100000111010000011111100000";
                        f_reg(342) <= "00011111101000000000000000000011";
                        f_reg(343) <= "00100000000111010000000000111100";
                        f_reg(344) <= "00010000000000000000000000000010";
                        f_reg(345) <= "00100000000111010000000000000000";
                        f_reg(346) <= "00010101000101100000000000110101";
                        f_reg(347) <= "10101111101010000000011110000100";
                        f_reg(348) <= "10001100000111010000011111100000";
                        f_reg(349) <= "00011111101000000000000000000011";
                        f_reg(350) <= "00100000000111010000000000111100";
                        f_reg(351) <= "00010000000000000000000000000010";
                        f_reg(352) <= "00100000000111010000000000000000";
                        f_reg(353) <= "00010101001101110000000000101110";
                        f_reg(354) <= "10101111101010010000011110001000";
                        f_reg(355) <= "10001100000111010000011111100000";
                        f_reg(356) <= "00011111101000000000000000000011";
                        f_reg(357) <= "00100000000111010000000000111100";
                        f_reg(358) <= "00010000000000000000000000000010";
                        f_reg(359) <= "00100000000111010000000000000000";
                        f_reg(360) <= "00010101010110000000000000100111";
                        f_reg(361) <= "10101111101010100000011110001100";
                        f_reg(362) <= "10001100000111010000011111100000";
                        f_reg(363) <= "00011111101000000000000000000011";
                        f_reg(364) <= "00100000000111010000000000111100";
                        f_reg(365) <= "00010000000000000000000000000010";
                        f_reg(366) <= "00100000000111010000000000000000";
                        f_reg(367) <= "00010101011110010000000000100000";
                        f_reg(368) <= "10101111101010110000011110010000";
                        f_reg(369) <= "10001100000111010000011111100000";
                        f_reg(370) <= "00011111101000000000000000000011";
                        f_reg(371) <= "00100000000111010000000000111100";
                        f_reg(372) <= "00010000000000000000000000000010";
                        f_reg(373) <= "00100000000111010000000000000000";
                        f_reg(374) <= "00010101100110100000000000011001";
                        f_reg(375) <= "10101111101011000000011110010100";
                        f_reg(376) <= "10001100000111010000011111100000";
                        f_reg(377) <= "00011111101000000000000000000011";
                        f_reg(378) <= "00100000000111010000000000111100";
                        f_reg(379) <= "00010000000000000000000000000010";
                        f_reg(380) <= "00100000000111010000000000000000";
                        f_reg(381) <= "00010101101110110000000000010010";
                        f_reg(382) <= "10101111101011010000011110011000";
                        f_reg(383) <= "10001100000111010000011111100000";
                        f_reg(384) <= "00011111101000000000000000000011";
                        f_reg(385) <= "00100000000111010000000000111100";
                        f_reg(386) <= "00010000000000000000000000000010";
                        f_reg(387) <= "00100000000111010000000000000000";
                        f_reg(388) <= "00010101110111000000000000001011";
                        f_reg(389) <= "10101111101011100000011110011100";
                        f_reg(390) <= "10001100000111010000011111100000";
                        f_reg(391) <= "00011111101000000000000000000011";
                        f_reg(392) <= "00100000000111010000000000111100";
                        f_reg(393) <= "00010000000000000000000000000010";
                        f_reg(394) <= "00100000000111010000000000000000";
                        f_reg(395) <= "00010111110111110000000000000100";
                        f_reg(396) <= "10101111101111100000011110100000";
                        f_reg(397) <= "10101100000111010000011111100000";
                        f_reg(398) <= "00010000000000001111111101111110";
                        f_reg(399) <= "10001100000111010000011111100000";
                        f_reg(400) <= "10001111101000010000011101101000";
                        f_reg(401) <= "10001100000111010000011111100000";
                        f_reg(402) <= "10001111101011110000011101101000";
                        f_reg(403) <= "00010100001011111111111111111100";
                        f_reg(404) <= "10001100000111010000011111100000";
                        f_reg(405) <= "10001111101000100000011101101100";
                        f_reg(406) <= "10001100000111010000011111100000";
                        f_reg(407) <= "10001111101100000000011101101100";
                        f_reg(408) <= "00010100010100001111111111111100";
                        f_reg(409) <= "10001100000111010000011111100000";
                        f_reg(410) <= "10001111101000110000011101110000";
                        f_reg(411) <= "10001100000111010000011111100000";
                        f_reg(412) <= "10001111101100010000011101110000";
                        f_reg(413) <= "00010100011100011111111111111100";
                        f_reg(414) <= "10001100000111010000011111100000";
                        f_reg(415) <= "10001111101001000000011101110100";
                        f_reg(416) <= "10001100000111010000011111100000";
                        f_reg(417) <= "10001111101100100000011101110100";
                        f_reg(418) <= "00010100100100101111111111111100";
                        f_reg(419) <= "10001100000111010000011111100000";
                        f_reg(420) <= "10001111101001010000011101111000";
                        f_reg(421) <= "10001100000111010000011111100000";
                        f_reg(422) <= "10001111101100110000011101111000";
                        f_reg(423) <= "00010100101100111111111111111100";
                        f_reg(424) <= "10001100000111010000011111100000";
                        f_reg(425) <= "10001111101001100000011101111100";
                        f_reg(426) <= "10001100000111010000011111100000";
                        f_reg(427) <= "10001111101101000000011101111100";
                        f_reg(428) <= "00010100110101001111111111111100";
                        f_reg(429) <= "10001100000111010000011111100000";
                        f_reg(430) <= "10001111101001110000011110000000";
                        f_reg(431) <= "10001100000111010000011111100000";
                        f_reg(432) <= "10001111101101010000011110000000";
                        f_reg(433) <= "00010100111101011111111111111100";
                        f_reg(434) <= "10001100000111010000011111100000";
                        f_reg(435) <= "10001111101010000000011110000100";
                        f_reg(436) <= "10001100000111010000011111100000";
                        f_reg(437) <= "10001111101101100000011110000100";
                        f_reg(438) <= "00010101000101101111111111111100";
                        f_reg(439) <= "10001100000111010000011111100000";
                        f_reg(440) <= "10001111101010010000011110001000";
                        f_reg(441) <= "10001100000111010000011111100000";
                        f_reg(442) <= "10001111101101110000011110001000";
                        f_reg(443) <= "00010101001101111111111111111100";
                        f_reg(444) <= "10001100000111010000011111100000";
                        f_reg(445) <= "10001111101010100000011110001100";
                        f_reg(446) <= "10001100000111010000011111100000";
                        f_reg(447) <= "10001111101110000000011110001100";
                        f_reg(448) <= "00010101010110001111111111111100";
                        f_reg(449) <= "10001100000111010000011111100000";
                        f_reg(450) <= "10001111101010110000011110010000";
                        f_reg(451) <= "10001100000111010000011111100000";
                        f_reg(452) <= "10001111101110010000011110010000";
                        f_reg(453) <= "00010101011110011111111111111100";
                        f_reg(454) <= "10001100000111010000011111100000";
                        f_reg(455) <= "10001111101011000000011110010100";
                        f_reg(456) <= "10001100000111010000011111100000";
                        f_reg(457) <= "10001111101110100000011110010100";
                        f_reg(458) <= "00010101100110101111111111111100";
                        f_reg(459) <= "10001100000111010000011111100000";
                        f_reg(460) <= "10001111101011010000011110011000";
                        f_reg(461) <= "10001100000111010000011111100000";
                        f_reg(462) <= "10001111101110110000011110011000";
                        f_reg(463) <= "00010101101110111111111111111100";
                        f_reg(464) <= "10001100000111010000011111100000";
                        f_reg(465) <= "10001111101011100000011110011100";
                        f_reg(466) <= "10001100000111010000011111100000";
                        f_reg(467) <= "10001111101111000000011110011100";
                        f_reg(468) <= "00010101110111001111111111111100";
                        f_reg(469) <= "10001100000111010000011111100000";
                        f_reg(470) <= "10001111101111100000011110100000";
                        f_reg(471) <= "10001100000111010000011111100000";
                        f_reg(472) <= "10001111101111110000011110100000";
                        f_reg(473) <= "00010111110111111111111111111100";
                        f_reg(474) <= "00010000000000001111111100110010";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000001111100111";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 4821
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SUB R2 R1 R1
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SLTI R3 R1 10399
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- ADD R4 R1 R1
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SRA R5 R2 1
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- SUBU R6 R5 R3
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- OR R7 R2 R2
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- SRA R8 R0 7
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- SW R8 R0 1088
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- SW R1 R0 1092
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- SRLV R9 R4 R4
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- SLTU R10 R7 R7
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- NOR R11 R6 R10
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- SW R8 R0 1096
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- SLLV R12 R1 R8
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- NOP
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SLTU R13 R12 R11
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- SRL R14 R8 6
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SW R1 R0 1100
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- SLTU R5 R9 R5
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- SUBU R15 R1 R6
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- AND R16 R4 R3
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- SLTI R17 R14 -30419
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- NOR R18 R4 R6
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- SLTIU R19 R8 18434
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- AND R20 R13 R1
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- SW R12 R0 1104
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- SRLV R21 R1 R0
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- ADDU R22 R18 R14
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- SLT R23 R5 R15
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- ADDU R24 R11 R10
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- SW R10 R0 1108
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- NOP
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- OR R25 R19 R18
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- SRA R26 R9 16
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- SW R25 R0 1112
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- SUB R6 R6 R4
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- ADDIU R27 R23 -11017
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- NOR R5 R5 R13
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- SRA R28 R25 16
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SLTIU R29 R11 5709
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- SLTU R30 R27 R16
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- ADD R2 R24 R18
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- AND R7 R20 R0
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- SW R7 R0 1116
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- ANDI R3 R21 -32648
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- SUBU R12 R2 R30
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- SUB R1 R26 R28
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SLTU R14 R6 R30
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- OR R15 R2 R8
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- ADDIU R10 R25 -32452
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- XORI R9 R5 -16051
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SW R17 R0 1120
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- SLTIU R4 R14 28127
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SW R15 R0 1124
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- SW R10 R0 1128
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- SLLV R23 R9 R30
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SLT R13 R3 R29
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- XOR R11 R1 R4
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- NOR R27 R6 R14
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- NOP
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- SW R27 R0 1132
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- SW R13 R0 1136
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- AND R16 R23 R0
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- SUB R24 R19 R12
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- ADD R18 R22 R11
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- NOP
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- ORI R20 R16 28741
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- NOP
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- SLTU R7 R20 R24
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SW R7 R0 1140
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- SLL R18 R18 15
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- NOP
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- SW R18 R0 1144
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- ADDI R31 R31 -1
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- BGTZ R31 -75
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- BEQ R0 R0 461
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- LUI R30 999
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- LUI R31 999
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- SRL R30 R30 16
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SRL R31 R31 16
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- LUI R1 4821
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- LUI R15 4821
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- SUB R2 R1 R1
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SUB R16 R15 R15
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- SLTI R3 R1 10399
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- SLTI R17 R15 10399
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- ADD R4 R1 R1
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- ADD R18 R15 R15
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- SRA R5 R2 1
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- SRA R19 R16 1
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- SUBU R6 R5 R3
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- SUBU R20 R19 R17
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- OR R7 R2 R2
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- OR R21 R16 R16
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SRA R8 R0 7
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- SRA R22 R0 7
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- BNE R8 R22 299
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- SW R8 R0 1088
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- BNE R1 R15 297
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SW R1 R0 1092
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- SRLV R9 R4 R4
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- SRLV R23 R18 R18
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- SLTU R10 R7 R7
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- SLTU R24 R21 R21
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- NOR R11 R6 R10
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- NOR R25 R20 R24
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- BNE R8 R22 289
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- SW R8 R0 1096
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- SLLV R12 R1 R8
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- SLLV R26 R15 R22
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- NOP
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- NOP
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- SLTU R13 R12 R11
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- SLTU R27 R26 R25
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- SRL R14 R8 6
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- SRL R28 R22 6
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- BNE R1 R15 279
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- SW R1 R0 1100
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- SLTU R5 R9 R5
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- SLTU R19 R23 R19
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SUBU R2 R1 R6
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- SUBU R16 R15 R20
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- AND R7 R4 R3
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- AND R21 R18 R17
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SLTI R3 R14 -30419
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- SLTI R17 R28 -30419
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- BNE R3 R17 269
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- SW R3 R0 1148
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- NOR R3 R4 R6
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- NOR R17 R18 R20
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- BNE R3 R17 265
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- SW R3 R0 1152
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- SLTIU R3 R8 18434
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- SLTIU R17 R22 18434
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- BNE R3 R17 261
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- SW R3 R0 1156
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- AND R3 R13 R1
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- AND R17 R27 R15
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- BNE R12 R26 257
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- SW R12 R0 1104
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- SRLV R12 R1 R0
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- SRLV R26 R15 R0
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- LW R1 R0 1152
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- LW R15 R0 1152
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- BNE R1 R15 -2
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- BNE R8 R22 250
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- SW R8 R0 1152
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- ADDU R8 R1 R14
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- ADDU R22 R15 R28
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- SLT R14 R5 R2
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- SLT R28 R19 R16
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- ADDU R2 R11 R10
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- ADDU R16 R25 R24
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- BNE R10 R24 242
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- SW R10 R0 1108
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- NOP
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- NOP
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- LW R10 R0 1156
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- LW R24 R0 1156
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- BNE R10 R24 -2
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- BNE R8 R22 235
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- SW R8 R0 1156
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- OR R8 R10 R1
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- OR R22 R24 R15
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- BNE R10 R24 231
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- SW R10 R0 1160
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- SRA R10 R9 16
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- SRA R24 R23 16
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- BNE R8 R22 227
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- SW R8 R0 1112
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- SUB R6 R6 R4
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- SUB R20 R20 R18
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- ADDIU R9 R14 -11017
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- ADDIU R23 R28 -11017
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- NOR R5 R5 R13
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- NOR R19 R19 R27
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- SRA R4 R8 16
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- SRA R18 R22 16
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SLTIU R14 R11 5709
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- SLTIU R28 R25 5709
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- SLTU R13 R9 R7
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- SLTU R27 R23 R21
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- ADD R11 R2 R1
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- ADD R25 R16 R15
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- AND R9 R3 R0
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- AND R23 R17 R0
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- BNE R9 R23 209
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- SW R9 R0 1116
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- ANDI R7 R12 -32648
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- ANDI R21 R26 -32648
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- SUBU R2 R11 R13
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- SUBU R16 R25 R27
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- SUB R1 R10 R4
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- SUB R15 R24 R18
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- SLTU R3 R6 R13
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- SLTU R17 R20 R27
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- LW R9 R0 1152
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- LW R23 R0 1152
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- BNE R9 R23 -2
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- OR R12 R11 R9
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- OR R26 R25 R23
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- ADDIU R10 R8 -32452
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- ADDIU R24 R22 -32452
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- XORI R4 R5 -16051
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- XORI R18 R19 -16051
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- LW R11 R0 1148
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- LW R25 R0 1148
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- BNE R11 R25 -2
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- BNE R11 R25 187
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- SW R11 R0 1120
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- SLTIU R9 R3 28127
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- SLTIU R23 R17 28127
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- BNE R12 R26 183
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- SW R12 R0 1124
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- BNE R10 R24 181
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- SW R10 R0 1128
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- SLLV R8 R4 R13
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- SLLV R22 R18 R27
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- SLT R5 R7 R14
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- SLT R19 R21 R28
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- XOR R11 R1 R9
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- XOR R25 R15 R23
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- NOR R12 R6 R3
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- NOR R26 R20 R17
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- NOP
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- NOP
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- BNE R12 R26 169
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- SW R12 R0 1132
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- BNE R5 R19 167
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- SW R5 R0 1136
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- AND R10 R8 R0
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- AND R24 R22 R0
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- LW R4 R0 1160
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- LW R18 R0 1160
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- BNE R4 R18 -2
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- SUB R13 R4 R2
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- SUB R27 R18 R16
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- LW R7 R0 1156
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- LW R21 R0 1156
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- BNE R7 R21 -2
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- ADD R14 R7 R11
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- ADD R28 R21 R25
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- NOP
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- NOP
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- ORI R1 R10 28741
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- ORI R15 R24 28741
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- NOP
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- NOP
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- SLTU R9 R1 R13
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- SLTU R23 R15 R27
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- BNE R9 R23 145
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- SW R9 R0 1140
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- SLL R14 R14 15
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- SLL R28 R28 15
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- NOP
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- NOP
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- BNE R14 R28 139
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- SW R14 R0 1144
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- ADDI R29 R30 -250
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- BEQ R29 R0 29
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- ADDI R29 R30 -500
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- BEQ R29 R0 27
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- ADDI R29 R30 -750
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- BEQ R29 R0 25
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- ADDI R30 R30 -1
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- ADDI R31 R31 -1
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- BNE R30 R31 129
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- BGTZ R31 -187
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- BEQ R0 R0 268
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- NOP
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- NOP
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- NOP
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- NOP
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- NOP
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- NOP
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- NOP
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- NOP
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- NOP
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- NOP
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- NOP
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- NOP
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- NOP
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- NOP
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- NOP
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- NOP
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- NOP
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- NOP
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- NOP
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- LW R29 R0 2016
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- BGTZ R29 3
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- ADDI R29 R0 60
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- BEQ R0 R0 2
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- ADDI R29 R0 0
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- BNE R1 R15 102
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- SW R1 R29 1896
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- LW R29 R0 2016
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- BGTZ R29 3
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- ADDI R29 R0 60
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- BEQ R0 R0 2
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- ADDI R29 R0 0
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- BNE R2 R16 95
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- SW R2 R29 1900
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- LW R29 R0 2016
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- BGTZ R29 3
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- ADDI R29 R0 60
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- BEQ R0 R0 2
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- ADDI R29 R0 0
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- BNE R3 R17 88
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- SW R3 R29 1904
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- LW R29 R0 2016
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- BGTZ R29 3
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- ADDI R29 R0 60
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- BEQ R0 R0 2
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- ADDI R29 R0 0
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- BNE R4 R18 81
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- SW R4 R29 1908
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- LW R29 R0 2016
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- BGTZ R29 3
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- ADDI R29 R0 60
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- BEQ R0 R0 2
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- ADDI R29 R0 0
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- BNE R5 R19 74
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- SW R5 R29 1912
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- LW R29 R0 2016
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- BGTZ R29 3
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- ADDI R29 R0 60
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- BEQ R0 R0 2
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- ADDI R29 R0 0
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- BNE R6 R20 67
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- SW R6 R29 1916
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- LW R29 R0 2016
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- BGTZ R29 3
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- ADDI R29 R0 60
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- BEQ R0 R0 2
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- ADDI R29 R0 0
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- BNE R7 R21 60
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- SW R7 R29 1920
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- LW R29 R0 2016
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- BGTZ R29 3
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- ADDI R29 R0 60
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- BEQ R0 R0 2
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- ADDI R29 R0 0
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- BNE R8 R22 53
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- SW R8 R29 1924
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- LW R29 R0 2016
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- BGTZ R29 3
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- ADDI R29 R0 60
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- BEQ R0 R0 2
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- ADDI R29 R0 0
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- BNE R9 R23 46
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- SW R9 R29 1928
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- LW R29 R0 2016
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- BGTZ R29 3
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- ADDI R29 R0 60
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- BEQ R0 R0 2
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- ADDI R29 R0 0
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- BNE R10 R24 39
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- SW R10 R29 1932
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- LW R29 R0 2016
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- BGTZ R29 3
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- ADDI R29 R0 60
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- BEQ R0 R0 2
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- ADDI R29 R0 0
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- BNE R11 R25 32
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- SW R11 R29 1936
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- LW R29 R0 2016
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- BGTZ R29 3
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- ADDI R29 R0 60
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- BEQ R0 R0 2
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- ADDI R29 R0 0
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- BNE R12 R26 25
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- SW R12 R29 1940
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- LW R29 R0 2016
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- BGTZ R29 3
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- ADDI R29 R0 60
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- BEQ R0 R0 2
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- ADDI R29 R0 0
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- BNE R13 R27 18
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- SW R13 R29 1944
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- LW R29 R0 2016
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- BGTZ R29 3
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- ADDI R29 R0 60
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- BEQ R0 R0 2
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- ADDI R29 R0 0
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- BNE R14 R28 11
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- SW R14 R29 1948
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- LW R29 R0 2016
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- BGTZ R29 3
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- ADDI R29 R0 60
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- BEQ R0 R0 2
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- ADDI R29 R0 0
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- BNE R30 R31 4
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- SW R30 R29 1952
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- SW R29 R0 2016
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- BEQ R0 R0 -130
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- LW R29 R0 2016
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- LW R1 R29 1896
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- LW R29 R0 2016
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- LW R15 R29 1896
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- BNE R1 R15 -4
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- LW R29 R0 2016
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- LW R2 R29 1900
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- LW R29 R0 2016
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- LW R16 R29 1900
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- BNE R2 R16 -4
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- LW R29 R0 2016
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- LW R3 R29 1904
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- LW R29 R0 2016
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- LW R17 R29 1904
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- BNE R3 R17 -4
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- LW R29 R0 2016
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- LW R4 R29 1908
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- LW R29 R0 2016
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- LW R18 R29 1908
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- BNE R4 R18 -4
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- LW R29 R0 2016
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- LW R5 R29 1912
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- LW R29 R0 2016
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- LW R19 R29 1912
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- BNE R5 R19 -4
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- LW R29 R0 2016
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R6 R29 1916
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R29 R0 2016
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- LW R20 R29 1916
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- BNE R6 R20 -4
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- LW R29 R0 2016
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- LW R7 R29 1920
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- LW R29 R0 2016
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- LW R21 R29 1920
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- BNE R7 R21 -4
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- LW R29 R0 2016
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- LW R8 R29 1924
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- LW R29 R0 2016
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- LW R22 R29 1924
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- BNE R8 R22 -4
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- LW R29 R0 2016
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- LW R9 R29 1928
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- LW R29 R0 2016
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- LW R23 R29 1928
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- BNE R9 R23 -4
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- LW R29 R0 2016
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- LW R10 R29 1932
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- LW R29 R0 2016
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- LW R24 R29 1932
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- BNE R10 R24 -4
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- LW R29 R0 2016
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- LW R11 R29 1936
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- LW R29 R0 2016
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- LW R25 R29 1936
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- BNE R11 R25 -4
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- LW R29 R0 2016
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- LW R12 R29 1940
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- LW R29 R0 2016
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- LW R26 R29 1940
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- BNE R12 R26 -4
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- LW R29 R0 2016
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- LW R13 R29 1944
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- LW R29 R0 2016
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- LW R27 R29 1944
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- BNE R13 R27 -4
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- LW R29 R0 2016
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- LW R14 R29 1948
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- LW R29 R0 2016
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- LW R28 R29 1948
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- BNE R14 R28 -4
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- LW R29 R0 2016
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- LW R30 R29 1952
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- LW R29 R0 2016
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- LW R31 R29 1952
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- BNE R30 R31 -4
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- BEQ R0 R0 -206
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- NOP
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- NOP
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- NOP
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- NOP
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- NOP
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- NOP
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- NOP
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- NOP
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- NOP
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- NOP
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- NOP
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- NOP
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- NOP
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- NOP
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- NOP
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- NOP
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- NOP
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- NOP
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- NOP
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- NOP
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- NOP
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- NOP
                        f_reg(496) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(497) =>
                        -- NOP
                        f_reg(497) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(498) =>
                        -- NOP
                        f_reg(498) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(499) =>
                        -- NOP
                        f_reg(499) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(500) =>
                        -- NOP
                        f_reg(500) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(501) =>
                        -- NOP
                        f_reg(501) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(502) =>
                        -- NOP
                        f_reg(502) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(503) =>
                        -- NOP
                        f_reg(503) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(504) =>
                        -- NOP
                        f_reg(504) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(505) =>
                        -- NOP
                        f_reg(505) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(506) =>
                        -- NOP
                        f_reg(506) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(507) =>
                        -- NOP
                        f_reg(507) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(508) =>
                        -- NOP
                        f_reg(508) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(509) =>
                        -- NOP
                        f_reg(509) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(510) =>
                        -- NOP
                        f_reg(510) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(511) =>
                        -- NOP
                        f_reg(511) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(512) =>
                        -- NOP
                        f_reg(512) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(513) =>
                        -- NOP
                        f_reg(513) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(514) =>
                        -- NOP
                        f_reg(514) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(515) =>
                        -- NOP
                        f_reg(515) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(516) =>
                        -- NOP
                        f_reg(516) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(517) =>
                        -- NOP
                        f_reg(517) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(518) =>
                        -- NOP
                        f_reg(518) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(519) =>
                        -- NOP
                        f_reg(519) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(520) =>
                        -- NOP
                        f_reg(520) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(521) =>
                        -- NOP
                        f_reg(521) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(522) =>
                        -- NOP
                        f_reg(522) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(523) =>
                        -- NOP
                        f_reg(523) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(524) =>
                        -- NOP
                        f_reg(524) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(525) =>
                        -- NOP
                        f_reg(525) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(526) =>
                        -- NOP
                        f_reg(526) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(527) =>
                        -- NOP
                        f_reg(527) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(528) =>
                        -- NOP
                        f_reg(528) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(529) =>
                        -- NOP
                        f_reg(529) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(530) =>
                        -- NOP
                        f_reg(530) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(531) =>
                        -- NOP
                        f_reg(531) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(532) =>
                        -- NOP
                        f_reg(532) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(533) =>
                        -- NOP
                        f_reg(533) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(534) =>
                        -- NOP
                        f_reg(534) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(535) =>
                        -- NOP
                        f_reg(535) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(536) =>
                        -- NOP
                        f_reg(536) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(537) =>
                        -- NOP
                        f_reg(537) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(538) =>
                        -- NOP
                        f_reg(538) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(539) =>
                        -- NOP
                        f_reg(539) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(540) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010001001011010101";
                        f_reg(4) <= "00000000001000010001000000100010";
                        f_reg(5) <= "00101000001000110010100010011111";
                        f_reg(6) <= "00000000001000010010000000100000";
                        f_reg(7) <= "00000000000000100010100001000011";
                        f_reg(8) <= "00000000101000110011000000100011";
                        f_reg(9) <= "00000000010000100011100000100101";
                        f_reg(10) <= "00000000000000000100000111000011";
                        f_reg(11) <= "10101100000010000000010001000000";
                        f_reg(12) <= "10101100000000010000010001000100";
                        f_reg(13) <= "00000000100001000100100000000110";
                        f_reg(14) <= "00000000111001110101000000101011";
                        f_reg(15) <= "00000000110010100101100000100111";
                        f_reg(16) <= "10101100000010000000010001001000";
                        f_reg(17) <= "00000001000000010110000000000100";
                        f_reg(18) <= "00000000000000000000000000000000";
                        f_reg(19) <= "00000001100010110110100000101011";
                        f_reg(20) <= "00000000000010000111000110000010";
                        f_reg(21) <= "10101100000000010000010001001100";
                        f_reg(22) <= "00000001001001010010100000101011";
                        f_reg(23) <= "00000000001001100111100000100011";
                        f_reg(24) <= "00000000100000111000000000100100";
                        f_reg(25) <= "00101001110100011000100100101101";
                        f_reg(26) <= "00000000100001101001000000100111";
                        f_reg(27) <= "00101101000100110100100000000010";
                        f_reg(28) <= "00000001101000011010000000100100";
                        f_reg(29) <= "10101100000011000000010001010000";
                        f_reg(30) <= "00000000000000011010100000000110";
                        f_reg(31) <= "00000010010011101011000000100001";
                        f_reg(32) <= "00000000101011111011100000101010";
                        f_reg(33) <= "00000001011010101100000000100001";
                        f_reg(34) <= "10101100000010100000010001010100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000010011100101100100000100101";
                        f_reg(37) <= "00000000000010011101010000000011";
                        f_reg(38) <= "10101100000110010000010001011000";
                        f_reg(39) <= "00000000110001000011000000100010";
                        f_reg(40) <= "00100110111110111101010011110111";
                        f_reg(41) <= "00000000101011010010100000100111";
                        f_reg(42) <= "00000000000110011110010000000011";
                        f_reg(43) <= "00101101011111010001011001001101";
                        f_reg(44) <= "00000011011100001111000000101011";
                        f_reg(45) <= "00000011000100100001000000100000";
                        f_reg(46) <= "00000010100000000011100000100100";
                        f_reg(47) <= "10101100000001110000010001011100";
                        f_reg(48) <= "00110010101000111000000001111000";
                        f_reg(49) <= "00000000010111100110000000100011";
                        f_reg(50) <= "00000011010111000000100000100010";
                        f_reg(51) <= "00000000110111100111000000101011";
                        f_reg(52) <= "00000000010010000111100000100101";
                        f_reg(53) <= "00100111001010101000000100111100";
                        f_reg(54) <= "00111000101010011100000101001101";
                        f_reg(55) <= "10101100000100010000010001100000";
                        f_reg(56) <= "00101101110001000110110111011111";
                        f_reg(57) <= "10101100000011110000010001100100";
                        f_reg(58) <= "10101100000010100000010001101000";
                        f_reg(59) <= "00000011110010011011100000000100";
                        f_reg(60) <= "00000000011111010110100000101010";
                        f_reg(61) <= "00000000001001000101100000100110";
                        f_reg(62) <= "00000000110011101101100000100111";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000110110000010001101100";
                        f_reg(65) <= "10101100000011010000010001110000";
                        f_reg(66) <= "00000010111000001000000000100100";
                        f_reg(67) <= "00000010011011001100000000100010";
                        f_reg(68) <= "00000010110010111001000000100000";
                        f_reg(69) <= "00000000000000000000000000000000";
                        f_reg(70) <= "00110110000101000111000001000101";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000010100110000011100000101011";
                        f_reg(73) <= "10101100000001110000010001110100";
                        f_reg(74) <= "00000000000100101001001111000000";
                        f_reg(75) <= "00000000000000000000000000000000";
                        f_reg(76) <= "10101100000100100000010001111000";
                        f_reg(77) <= "00100011111111111111111111111111";
                        f_reg(78) <= "00011111111000001111111110110101";
                        f_reg(79) <= "00010000000000000000000111001101";
                        f_reg(80) <= "00111100000111100000001111100111";
                        f_reg(81) <= "00111100000111110000001111100111";
                        f_reg(82) <= "00000000000111101111010000000010";
                        f_reg(83) <= "00000000000111111111110000000010";
                        f_reg(84) <= "00111100000000010001001011010101";
                        f_reg(85) <= "00111100000011110001001011010101";
                        f_reg(86) <= "00000000001000010001000000100010";
                        f_reg(87) <= "00000001111011111000000000100010";
                        f_reg(88) <= "00101000001000110010100010011111";
                        f_reg(89) <= "00101001111100010010100010011111";
                        f_reg(90) <= "00000000001000010010000000100000";
                        f_reg(91) <= "00000001111011111001000000100000";
                        f_reg(92) <= "00000000000000100010100001000011";
                        f_reg(93) <= "00000000000100001001100001000011";
                        f_reg(94) <= "00000000101000110011000000100011";
                        f_reg(95) <= "00000010011100011010000000100011";
                        f_reg(96) <= "00000000010000100011100000100101";
                        f_reg(97) <= "00000010000100001010100000100101";
                        f_reg(98) <= "00000000000000000100000111000011";
                        f_reg(99) <= "00000000000000001011000111000011";
                        f_reg(100) <= "00010101000101100000000100101011";
                        f_reg(101) <= "10101100000010000000010001000000";
                        f_reg(102) <= "00010100001011110000000100101001";
                        f_reg(103) <= "10101100000000010000010001000100";
                        f_reg(104) <= "00000000100001000100100000000110";
                        f_reg(105) <= "00000010010100101011100000000110";
                        f_reg(106) <= "00000000111001110101000000101011";
                        f_reg(107) <= "00000010101101011100000000101011";
                        f_reg(108) <= "00000000110010100101100000100111";
                        f_reg(109) <= "00000010100110001100100000100111";
                        f_reg(110) <= "00010101000101100000000100100001";
                        f_reg(111) <= "10101100000010000000010001001000";
                        f_reg(112) <= "00000001000000010110000000000100";
                        f_reg(113) <= "00000010110011111101000000000100";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00000000000000000000000000000000";
                        f_reg(116) <= "00000001100010110110100000101011";
                        f_reg(117) <= "00000011010110011101100000101011";
                        f_reg(118) <= "00000000000010000111000110000010";
                        f_reg(119) <= "00000000000101101110000110000010";
                        f_reg(120) <= "00010100001011110000000100010111";
                        f_reg(121) <= "10101100000000010000010001001100";
                        f_reg(122) <= "00000001001001010010100000101011";
                        f_reg(123) <= "00000010111100111001100000101011";
                        f_reg(124) <= "00000000001001100001000000100011";
                        f_reg(125) <= "00000001111101001000000000100011";
                        f_reg(126) <= "00000000100000110011100000100100";
                        f_reg(127) <= "00000010010100011010100000100100";
                        f_reg(128) <= "00101001110000111000100100101101";
                        f_reg(129) <= "00101011100100011000100100101101";
                        f_reg(130) <= "00010100011100010000000100001101";
                        f_reg(131) <= "10101100000000110000010001111100";
                        f_reg(132) <= "00000000100001100001100000100111";
                        f_reg(133) <= "00000010010101001000100000100111";
                        f_reg(134) <= "00010100011100010000000100001001";
                        f_reg(135) <= "10101100000000110000010010000000";
                        f_reg(136) <= "00101101000000110100100000000010";
                        f_reg(137) <= "00101110110100010100100000000010";
                        f_reg(138) <= "00010100011100010000000100000101";
                        f_reg(139) <= "10101100000000110000010010000100";
                        f_reg(140) <= "00000001101000010001100000100100";
                        f_reg(141) <= "00000011011011111000100000100100";
                        f_reg(142) <= "00010101100110100000000100000001";
                        f_reg(143) <= "10101100000011000000010001010000";
                        f_reg(144) <= "00000000000000010110000000000110";
                        f_reg(145) <= "00000000000011111101000000000110";
                        f_reg(146) <= "10001100000000010000010010000000";
                        f_reg(147) <= "10001100000011110000010010000000";
                        f_reg(148) <= "00010100001011111111111111111110";
                        f_reg(149) <= "00010101000101100000000011111010";
                        f_reg(150) <= "10101100000010000000010010000000";
                        f_reg(151) <= "00000000001011100100000000100001";
                        f_reg(152) <= "00000001111111001011000000100001";
                        f_reg(153) <= "00000000101000100111000000101010";
                        f_reg(154) <= "00000010011100001110000000101010";
                        f_reg(155) <= "00000001011010100001000000100001";
                        f_reg(156) <= "00000011001110001000000000100001";
                        f_reg(157) <= "00010101010110000000000011110010";
                        f_reg(158) <= "10101100000010100000010001010100";
                        f_reg(159) <= "00000000000000000000000000000000";
                        f_reg(160) <= "00000000000000000000000000000000";
                        f_reg(161) <= "10001100000010100000010010000100";
                        f_reg(162) <= "10001100000110000000010010000100";
                        f_reg(163) <= "00010101010110001111111111111110";
                        f_reg(164) <= "00010101000101100000000011101011";
                        f_reg(165) <= "10101100000010000000010010000100";
                        f_reg(166) <= "00000001010000010100000000100101";
                        f_reg(167) <= "00000011000011111011000000100101";
                        f_reg(168) <= "00010101010110000000000011100111";
                        f_reg(169) <= "10101100000010100000010010001000";
                        f_reg(170) <= "00000000000010010101010000000011";
                        f_reg(171) <= "00000000000101111100010000000011";
                        f_reg(172) <= "00010101000101100000000011100011";
                        f_reg(173) <= "10101100000010000000010001011000";
                        f_reg(174) <= "00000000110001000011000000100010";
                        f_reg(175) <= "00000010100100101010000000100010";
                        f_reg(176) <= "00100101110010011101010011110111";
                        f_reg(177) <= "00100111100101111101010011110111";
                        f_reg(178) <= "00000000101011010010100000100111";
                        f_reg(179) <= "00000010011110111001100000100111";
                        f_reg(180) <= "00000000000010000010010000000011";
                        f_reg(181) <= "00000000000101101001010000000011";
                        f_reg(182) <= "00101101011011100001011001001101";
                        f_reg(183) <= "00101111001111000001011001001101";
                        f_reg(184) <= "00000001001001110110100000101011";
                        f_reg(185) <= "00000010111101011101100000101011";
                        f_reg(186) <= "00000000010000010101100000100000";
                        f_reg(187) <= "00000010000011111100100000100000";
                        f_reg(188) <= "00000000011000000100100000100100";
                        f_reg(189) <= "00000010001000001011100000100100";
                        f_reg(190) <= "00010101001101110000000011010001";
                        f_reg(191) <= "10101100000010010000010001011100";
                        f_reg(192) <= "00110001100001111000000001111000";
                        f_reg(193) <= "00110011010101011000000001111000";
                        f_reg(194) <= "00000001011011010001000000100011";
                        f_reg(195) <= "00000011001110111000000000100011";
                        f_reg(196) <= "00000001010001000000100000100010";
                        f_reg(197) <= "00000011000100100111100000100010";
                        f_reg(198) <= "00000000110011010001100000101011";
                        f_reg(199) <= "00000010100110111000100000101011";
                        f_reg(200) <= "10001100000010010000010010000000";
                        f_reg(201) <= "10001100000101110000010010000000";
                        f_reg(202) <= "00010101001101111111111111111110";
                        f_reg(203) <= "00000001011010010110000000100101";
                        f_reg(204) <= "00000011001101111101000000100101";
                        f_reg(205) <= "00100101000010101000000100111100";
                        f_reg(206) <= "00100110110110001000000100111100";
                        f_reg(207) <= "00111000101001001100000101001101";
                        f_reg(208) <= "00111010011100101100000101001101";
                        f_reg(209) <= "10001100000010110000010001111100";
                        f_reg(210) <= "10001100000110010000010001111100";
                        f_reg(211) <= "00010101011110011111111111111110";
                        f_reg(212) <= "00010101011110010000000010111011";
                        f_reg(213) <= "10101100000010110000010001100000";
                        f_reg(214) <= "00101100011010010110110111011111";
                        f_reg(215) <= "00101110001101110110110111011111";
                        f_reg(216) <= "00010101100110100000000010110111";
                        f_reg(217) <= "10101100000011000000010001100100";
                        f_reg(218) <= "00010101010110000000000010110101";
                        f_reg(219) <= "10101100000010100000010001101000";
                        f_reg(220) <= "00000001101001000100000000000100";
                        f_reg(221) <= "00000011011100101011000000000100";
                        f_reg(222) <= "00000000111011100010100000101010";
                        f_reg(223) <= "00000010101111001001100000101010";
                        f_reg(224) <= "00000000001010010101100000100110";
                        f_reg(225) <= "00000001111101111100100000100110";
                        f_reg(226) <= "00000000110000110110000000100111";
                        f_reg(227) <= "00000010100100011101000000100111";
                        f_reg(228) <= "00000000000000000000000000000000";
                        f_reg(229) <= "00000000000000000000000000000000";
                        f_reg(230) <= "00010101100110100000000010101001";
                        f_reg(231) <= "10101100000011000000010001101100";
                        f_reg(232) <= "00010100101100110000000010100111";
                        f_reg(233) <= "10101100000001010000010001110000";
                        f_reg(234) <= "00000001000000000101000000100100";
                        f_reg(235) <= "00000010110000001100000000100100";
                        f_reg(236) <= "10001100000001000000010010001000";
                        f_reg(237) <= "10001100000100100000010010001000";
                        f_reg(238) <= "00010100100100101111111111111110";
                        f_reg(239) <= "00000000100000100110100000100010";
                        f_reg(240) <= "00000010010100001101100000100010";
                        f_reg(241) <= "10001100000001110000010010000100";
                        f_reg(242) <= "10001100000101010000010010000100";
                        f_reg(243) <= "00010100111101011111111111111110";
                        f_reg(244) <= "00000000111010110111000000100000";
                        f_reg(245) <= "00000010101110011110000000100000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00110101010000010111000001000101";
                        f_reg(249) <= "00110111000011110111000001000101";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00000000000000000000000000000000";
                        f_reg(252) <= "00000000001011010100100000101011";
                        f_reg(253) <= "00000001111110111011100000101011";
                        f_reg(254) <= "00010101001101110000000010010001";
                        f_reg(255) <= "10101100000010010000010001110100";
                        f_reg(256) <= "00000000000011100111001111000000";
                        f_reg(257) <= "00000000000111001110001111000000";
                        f_reg(258) <= "00000000000000000000000000000000";
                        f_reg(259) <= "00000000000000000000000000000000";
                        f_reg(260) <= "00010101110111000000000010001011";
                        f_reg(261) <= "10101100000011100000010001111000";
                        f_reg(262) <= "00100011110111011111111100000110";
                        f_reg(263) <= "00010011101000000000000000011101";
                        f_reg(264) <= "00100011110111011111111000001100";
                        f_reg(265) <= "00010011101000000000000000011011";
                        f_reg(266) <= "00100011110111011111110100010010";
                        f_reg(267) <= "00010011101000000000000000011001";
                        f_reg(268) <= "00100011110111101111111111111111";
                        f_reg(269) <= "00100011111111111111111111111111";
                        f_reg(270) <= "00010111110111110000000010000001";
                        f_reg(271) <= "00011111111000001111111101000101";
                        f_reg(272) <= "00010000000000000000000100001100";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "00000000000000000000000000000000";
                        f_reg(287) <= "00000000000000000000000000000000";
                        f_reg(288) <= "00000000000000000000000000000000";
                        f_reg(289) <= "00000000000000000000000000000000";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "10001100000111010000011111100000";
                        f_reg(293) <= "00011111101000000000000000000011";
                        f_reg(294) <= "00100000000111010000000000111100";
                        f_reg(295) <= "00010000000000000000000000000010";
                        f_reg(296) <= "00100000000111010000000000000000";
                        f_reg(297) <= "00010100001011110000000001100110";
                        f_reg(298) <= "10101111101000010000011101101000";
                        f_reg(299) <= "10001100000111010000011111100000";
                        f_reg(300) <= "00011111101000000000000000000011";
                        f_reg(301) <= "00100000000111010000000000111100";
                        f_reg(302) <= "00010000000000000000000000000010";
                        f_reg(303) <= "00100000000111010000000000000000";
                        f_reg(304) <= "00010100010100000000000001011111";
                        f_reg(305) <= "10101111101000100000011101101100";
                        f_reg(306) <= "10001100000111010000011111100000";
                        f_reg(307) <= "00011111101000000000000000000011";
                        f_reg(308) <= "00100000000111010000000000111100";
                        f_reg(309) <= "00010000000000000000000000000010";
                        f_reg(310) <= "00100000000111010000000000000000";
                        f_reg(311) <= "00010100011100010000000001011000";
                        f_reg(312) <= "10101111101000110000011101110000";
                        f_reg(313) <= "10001100000111010000011111100000";
                        f_reg(314) <= "00011111101000000000000000000011";
                        f_reg(315) <= "00100000000111010000000000111100";
                        f_reg(316) <= "00010000000000000000000000000010";
                        f_reg(317) <= "00100000000111010000000000000000";
                        f_reg(318) <= "00010100100100100000000001010001";
                        f_reg(319) <= "10101111101001000000011101110100";
                        f_reg(320) <= "10001100000111010000011111100000";
                        f_reg(321) <= "00011111101000000000000000000011";
                        f_reg(322) <= "00100000000111010000000000111100";
                        f_reg(323) <= "00010000000000000000000000000010";
                        f_reg(324) <= "00100000000111010000000000000000";
                        f_reg(325) <= "00010100101100110000000001001010";
                        f_reg(326) <= "10101111101001010000011101111000";
                        f_reg(327) <= "10001100000111010000011111100000";
                        f_reg(328) <= "00011111101000000000000000000011";
                        f_reg(329) <= "00100000000111010000000000111100";
                        f_reg(330) <= "00010000000000000000000000000010";
                        f_reg(331) <= "00100000000111010000000000000000";
                        f_reg(332) <= "00010100110101000000000001000011";
                        f_reg(333) <= "10101111101001100000011101111100";
                        f_reg(334) <= "10001100000111010000011111100000";
                        f_reg(335) <= "00011111101000000000000000000011";
                        f_reg(336) <= "00100000000111010000000000111100";
                        f_reg(337) <= "00010000000000000000000000000010";
                        f_reg(338) <= "00100000000111010000000000000000";
                        f_reg(339) <= "00010100111101010000000000111100";
                        f_reg(340) <= "10101111101001110000011110000000";
                        f_reg(341) <= "10001100000111010000011111100000";
                        f_reg(342) <= "00011111101000000000000000000011";
                        f_reg(343) <= "00100000000111010000000000111100";
                        f_reg(344) <= "00010000000000000000000000000010";
                        f_reg(345) <= "00100000000111010000000000000000";
                        f_reg(346) <= "00010101000101100000000000110101";
                        f_reg(347) <= "10101111101010000000011110000100";
                        f_reg(348) <= "10001100000111010000011111100000";
                        f_reg(349) <= "00011111101000000000000000000011";
                        f_reg(350) <= "00100000000111010000000000111100";
                        f_reg(351) <= "00010000000000000000000000000010";
                        f_reg(352) <= "00100000000111010000000000000000";
                        f_reg(353) <= "00010101001101110000000000101110";
                        f_reg(354) <= "10101111101010010000011110001000";
                        f_reg(355) <= "10001100000111010000011111100000";
                        f_reg(356) <= "00011111101000000000000000000011";
                        f_reg(357) <= "00100000000111010000000000111100";
                        f_reg(358) <= "00010000000000000000000000000010";
                        f_reg(359) <= "00100000000111010000000000000000";
                        f_reg(360) <= "00010101010110000000000000100111";
                        f_reg(361) <= "10101111101010100000011110001100";
                        f_reg(362) <= "10001100000111010000011111100000";
                        f_reg(363) <= "00011111101000000000000000000011";
                        f_reg(364) <= "00100000000111010000000000111100";
                        f_reg(365) <= "00010000000000000000000000000010";
                        f_reg(366) <= "00100000000111010000000000000000";
                        f_reg(367) <= "00010101011110010000000000100000";
                        f_reg(368) <= "10101111101010110000011110010000";
                        f_reg(369) <= "10001100000111010000011111100000";
                        f_reg(370) <= "00011111101000000000000000000011";
                        f_reg(371) <= "00100000000111010000000000111100";
                        f_reg(372) <= "00010000000000000000000000000010";
                        f_reg(373) <= "00100000000111010000000000000000";
                        f_reg(374) <= "00010101100110100000000000011001";
                        f_reg(375) <= "10101111101011000000011110010100";
                        f_reg(376) <= "10001100000111010000011111100000";
                        f_reg(377) <= "00011111101000000000000000000011";
                        f_reg(378) <= "00100000000111010000000000111100";
                        f_reg(379) <= "00010000000000000000000000000010";
                        f_reg(380) <= "00100000000111010000000000000000";
                        f_reg(381) <= "00010101101110110000000000010010";
                        f_reg(382) <= "10101111101011010000011110011000";
                        f_reg(383) <= "10001100000111010000011111100000";
                        f_reg(384) <= "00011111101000000000000000000011";
                        f_reg(385) <= "00100000000111010000000000111100";
                        f_reg(386) <= "00010000000000000000000000000010";
                        f_reg(387) <= "00100000000111010000000000000000";
                        f_reg(388) <= "00010101110111000000000000001011";
                        f_reg(389) <= "10101111101011100000011110011100";
                        f_reg(390) <= "10001100000111010000011111100000";
                        f_reg(391) <= "00011111101000000000000000000011";
                        f_reg(392) <= "00100000000111010000000000111100";
                        f_reg(393) <= "00010000000000000000000000000010";
                        f_reg(394) <= "00100000000111010000000000000000";
                        f_reg(395) <= "00010111110111110000000000000100";
                        f_reg(396) <= "10101111101111100000011110100000";
                        f_reg(397) <= "10101100000111010000011111100000";
                        f_reg(398) <= "00010000000000001111111101111110";
                        f_reg(399) <= "10001100000111010000011111100000";
                        f_reg(400) <= "10001111101000010000011101101000";
                        f_reg(401) <= "10001100000111010000011111100000";
                        f_reg(402) <= "10001111101011110000011101101000";
                        f_reg(403) <= "00010100001011111111111111111100";
                        f_reg(404) <= "10001100000111010000011111100000";
                        f_reg(405) <= "10001111101000100000011101101100";
                        f_reg(406) <= "10001100000111010000011111100000";
                        f_reg(407) <= "10001111101100000000011101101100";
                        f_reg(408) <= "00010100010100001111111111111100";
                        f_reg(409) <= "10001100000111010000011111100000";
                        f_reg(410) <= "10001111101000110000011101110000";
                        f_reg(411) <= "10001100000111010000011111100000";
                        f_reg(412) <= "10001111101100010000011101110000";
                        f_reg(413) <= "00010100011100011111111111111100";
                        f_reg(414) <= "10001100000111010000011111100000";
                        f_reg(415) <= "10001111101001000000011101110100";
                        f_reg(416) <= "10001100000111010000011111100000";
                        f_reg(417) <= "10001111101100100000011101110100";
                        f_reg(418) <= "00010100100100101111111111111100";
                        f_reg(419) <= "10001100000111010000011111100000";
                        f_reg(420) <= "10001111101001010000011101111000";
                        f_reg(421) <= "10001100000111010000011111100000";
                        f_reg(422) <= "10001111101100110000011101111000";
                        f_reg(423) <= "00010100101100111111111111111100";
                        f_reg(424) <= "10001100000111010000011111100000";
                        f_reg(425) <= "10001111101001100000011101111100";
                        f_reg(426) <= "10001100000111010000011111100000";
                        f_reg(427) <= "10001111101101000000011101111100";
                        f_reg(428) <= "00010100110101001111111111111100";
                        f_reg(429) <= "10001100000111010000011111100000";
                        f_reg(430) <= "10001111101001110000011110000000";
                        f_reg(431) <= "10001100000111010000011111100000";
                        f_reg(432) <= "10001111101101010000011110000000";
                        f_reg(433) <= "00010100111101011111111111111100";
                        f_reg(434) <= "10001100000111010000011111100000";
                        f_reg(435) <= "10001111101010000000011110000100";
                        f_reg(436) <= "10001100000111010000011111100000";
                        f_reg(437) <= "10001111101101100000011110000100";
                        f_reg(438) <= "00010101000101101111111111111100";
                        f_reg(439) <= "10001100000111010000011111100000";
                        f_reg(440) <= "10001111101010010000011110001000";
                        f_reg(441) <= "10001100000111010000011111100000";
                        f_reg(442) <= "10001111101101110000011110001000";
                        f_reg(443) <= "00010101001101111111111111111100";
                        f_reg(444) <= "10001100000111010000011111100000";
                        f_reg(445) <= "10001111101010100000011110001100";
                        f_reg(446) <= "10001100000111010000011111100000";
                        f_reg(447) <= "10001111101110000000011110001100";
                        f_reg(448) <= "00010101010110001111111111111100";
                        f_reg(449) <= "10001100000111010000011111100000";
                        f_reg(450) <= "10001111101010110000011110010000";
                        f_reg(451) <= "10001100000111010000011111100000";
                        f_reg(452) <= "10001111101110010000011110010000";
                        f_reg(453) <= "00010101011110011111111111111100";
                        f_reg(454) <= "10001100000111010000011111100000";
                        f_reg(455) <= "10001111101011000000011110010100";
                        f_reg(456) <= "10001100000111010000011111100000";
                        f_reg(457) <= "10001111101110100000011110010100";
                        f_reg(458) <= "00010101100110101111111111111100";
                        f_reg(459) <= "10001100000111010000011111100000";
                        f_reg(460) <= "10001111101011010000011110011000";
                        f_reg(461) <= "10001100000111010000011111100000";
                        f_reg(462) <= "10001111101110110000011110011000";
                        f_reg(463) <= "00010101101110111111111111111100";
                        f_reg(464) <= "10001100000111010000011111100000";
                        f_reg(465) <= "10001111101011100000011110011100";
                        f_reg(466) <= "10001100000111010000011111100000";
                        f_reg(467) <= "10001111101111000000011110011100";
                        f_reg(468) <= "00010101110111001111111111111100";
                        f_reg(469) <= "10001100000111010000011111100000";
                        f_reg(470) <= "10001111101111100000011110100000";
                        f_reg(471) <= "10001100000111010000011111100000";
                        f_reg(472) <= "10001111101111110000011110100000";
                        f_reg(473) <= "00010111110111111111111111111100";
                        f_reg(474) <= "00010000000000001111111100110010";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000001111100111";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010001001011010101";
                        f_reg(4) <= "00000000001000010001000000100010";
                        f_reg(5) <= "00101000001000110010100010011111";
                        f_reg(6) <= "00000000001000010010000000100000";
                        f_reg(7) <= "00000000000000100010100001000011";
                        f_reg(8) <= "00000000101000110011000000100011";
                        f_reg(9) <= "00000000010000100011100000100101";
                        f_reg(10) <= "00000000000000000100000111000011";
                        f_reg(11) <= "10101100000010000000010001000000";
                        f_reg(12) <= "10101100000000010000010001000100";
                        f_reg(13) <= "00000000100001000100100000000110";
                        f_reg(14) <= "00000000111001110101000000101011";
                        f_reg(15) <= "00000000110010100101100000100111";
                        f_reg(16) <= "10101100000010000000010001001000";
                        f_reg(17) <= "00000001000000010110000000000100";
                        f_reg(18) <= "00000000000000000000000000000000";
                        f_reg(19) <= "00000001100010110110100000101011";
                        f_reg(20) <= "00000000000010000111000110000010";
                        f_reg(21) <= "10101100000000010000010001001100";
                        f_reg(22) <= "00000001001001010010100000101011";
                        f_reg(23) <= "00000000001001100111100000100011";
                        f_reg(24) <= "00000000100000111000000000100100";
                        f_reg(25) <= "00101001110100011000100100101101";
                        f_reg(26) <= "00000000100001101001000000100111";
                        f_reg(27) <= "00101101000100110100100000000010";
                        f_reg(28) <= "00000001101000011010000000100100";
                        f_reg(29) <= "10101100000011000000010001010000";
                        f_reg(30) <= "00000000000000011010100000000110";
                        f_reg(31) <= "00000010010011101011000000100001";
                        f_reg(32) <= "00000000101011111011100000101010";
                        f_reg(33) <= "00000001011010101100000000100001";
                        f_reg(34) <= "10101100000010100000010001010100";
                        f_reg(35) <= "00000000000000000000000000000000";
                        f_reg(36) <= "00000010011100101100100000100101";
                        f_reg(37) <= "00000000000010011101010000000011";
                        f_reg(38) <= "10101100000110010000010001011000";
                        f_reg(39) <= "00000000110001000011000000100010";
                        f_reg(40) <= "00100110111110111101010011110111";
                        f_reg(41) <= "00000000101011010010100000100111";
                        f_reg(42) <= "00000000000110011110010000000011";
                        f_reg(43) <= "00101101011111010001011001001101";
                        f_reg(44) <= "00000011011100001111000000101011";
                        f_reg(45) <= "00000011000100100001000000100000";
                        f_reg(46) <= "00000010100000000011100000100100";
                        f_reg(47) <= "10101100000001110000010001011100";
                        f_reg(48) <= "00110010101000111000000001111000";
                        f_reg(49) <= "00000000010111100110000000100011";
                        f_reg(50) <= "00000011010111000000100000100010";
                        f_reg(51) <= "00000000110111100111000000101011";
                        f_reg(52) <= "00000000010010000111100000100101";
                        f_reg(53) <= "00100111001010101000000100111100";
                        f_reg(54) <= "00111000101010011100000101001101";
                        f_reg(55) <= "10101100000100010000010001100000";
                        f_reg(56) <= "00101101110001000110110111011111";
                        f_reg(57) <= "10101100000011110000010001100100";
                        f_reg(58) <= "10101100000010100000010001101000";
                        f_reg(59) <= "00000011110010011011100000000100";
                        f_reg(60) <= "00000000011111010110100000101010";
                        f_reg(61) <= "00000000001001000101100000100110";
                        f_reg(62) <= "00000000110011101101100000100111";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000110110000010001101100";
                        f_reg(65) <= "10101100000011010000010001110000";
                        f_reg(66) <= "00000010111000001000000000100100";
                        f_reg(67) <= "00000010011011001100000000100010";
                        f_reg(68) <= "00000010110010111001000000100000";
                        f_reg(69) <= "00000000000000000000000000000000";
                        f_reg(70) <= "00110110000101000111000001000101";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000010100110000011100000101011";
                        f_reg(73) <= "10101100000001110000010001110100";
                        f_reg(74) <= "00000000000100101001001111000000";
                        f_reg(75) <= "00000000000000000000000000000000";
                        f_reg(76) <= "10101100000100100000010001111000";
                        f_reg(77) <= "00100011111111111111111111111111";
                        f_reg(78) <= "00011111111000001111111110110101";
                        f_reg(79) <= "00010000000000000000000111001101";
                        f_reg(80) <= "00111100000111100000001111100111";
                        f_reg(81) <= "00111100000111110000001111100111";
                        f_reg(82) <= "00000000000111101111010000000010";
                        f_reg(83) <= "00000000000111111111110000000010";
                        f_reg(84) <= "00111100000000010001001011010101";
                        f_reg(85) <= "00111100000011110001001011010101";
                        f_reg(86) <= "00000000001000010001000000100010";
                        f_reg(87) <= "00000001111011111000000000100010";
                        f_reg(88) <= "00101000001000110010100010011111";
                        f_reg(89) <= "00101001111100010010100010011111";
                        f_reg(90) <= "00000000001000010010000000100000";
                        f_reg(91) <= "00000001111011111001000000100000";
                        f_reg(92) <= "00000000000000100010100001000011";
                        f_reg(93) <= "00000000000100001001100001000011";
                        f_reg(94) <= "00000000101000110011000000100011";
                        f_reg(95) <= "00000010011100011010000000100011";
                        f_reg(96) <= "00000000010000100011100000100101";
                        f_reg(97) <= "00000010000100001010100000100101";
                        f_reg(98) <= "00000000000000000100000111000011";
                        f_reg(99) <= "00000000000000001011000111000011";
                        f_reg(100) <= "00010101000101100000000100101011";
                        f_reg(101) <= "10101100000010000000010001000000";
                        f_reg(102) <= "00010100001011110000000100101001";
                        f_reg(103) <= "10101100000000010000010001000100";
                        f_reg(104) <= "00000000100001000100100000000110";
                        f_reg(105) <= "00000010010100101011100000000110";
                        f_reg(106) <= "00000000111001110101000000101011";
                        f_reg(107) <= "00000010101101011100000000101011";
                        f_reg(108) <= "00000000110010100101100000100111";
                        f_reg(109) <= "00000010100110001100100000100111";
                        f_reg(110) <= "00010101000101100000000100100001";
                        f_reg(111) <= "10101100000010000000010001001000";
                        f_reg(112) <= "00000001000000010110000000000100";
                        f_reg(113) <= "00000010110011111101000000000100";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00000000000000000000000000000000";
                        f_reg(116) <= "00000001100010110110100000101011";
                        f_reg(117) <= "00000011010110011101100000101011";
                        f_reg(118) <= "00000000000010000111000110000010";
                        f_reg(119) <= "00000000000101101110000110000010";
                        f_reg(120) <= "00010100001011110000000100010111";
                        f_reg(121) <= "10101100000000010000010001001100";
                        f_reg(122) <= "00000001001001010010100000101011";
                        f_reg(123) <= "00000010111100111001100000101011";
                        f_reg(124) <= "00000000001001100001000000100011";
                        f_reg(125) <= "00000001111101001000000000100011";
                        f_reg(126) <= "00000000100000110011100000100100";
                        f_reg(127) <= "00000010010100011010100000100100";
                        f_reg(128) <= "00101001110000111000100100101101";
                        f_reg(129) <= "00101011100100011000100100101101";
                        f_reg(130) <= "00010100011100010000000100001101";
                        f_reg(131) <= "10101100000000110000010001111100";
                        f_reg(132) <= "00000000100001100001100000100111";
                        f_reg(133) <= "00000010010101001000100000100111";
                        f_reg(134) <= "00010100011100010000000100001001";
                        f_reg(135) <= "10101100000000110000010010000000";
                        f_reg(136) <= "00101101000000110100100000000010";
                        f_reg(137) <= "00101110110100010100100000000010";
                        f_reg(138) <= "00010100011100010000000100000101";
                        f_reg(139) <= "10101100000000110000010010000100";
                        f_reg(140) <= "00000001101000010001100000100100";
                        f_reg(141) <= "00000011011011111000100000100100";
                        f_reg(142) <= "00010101100110100000000100000001";
                        f_reg(143) <= "10101100000011000000010001010000";
                        f_reg(144) <= "00000000000000010110000000000110";
                        f_reg(145) <= "00000000000011111101000000000110";
                        f_reg(146) <= "10001100000000010000010010000000";
                        f_reg(147) <= "10001100000011110000010010000000";
                        f_reg(148) <= "00010100001011111111111111111110";
                        f_reg(149) <= "00010101000101100000000011111010";
                        f_reg(150) <= "10101100000010000000010010000000";
                        f_reg(151) <= "00000000001011100100000000100001";
                        f_reg(152) <= "00000001111111001011000000100001";
                        f_reg(153) <= "00000000101000100111000000101010";
                        f_reg(154) <= "00000010011100001110000000101010";
                        f_reg(155) <= "00000001011010100001000000100001";
                        f_reg(156) <= "00000011001110001000000000100001";
                        f_reg(157) <= "00010101010110000000000011110010";
                        f_reg(158) <= "10101100000010100000010001010100";
                        f_reg(159) <= "00000000000000000000000000000000";
                        f_reg(160) <= "00000000000000000000000000000000";
                        f_reg(161) <= "10001100000010100000010010000100";
                        f_reg(162) <= "10001100000110000000010010000100";
                        f_reg(163) <= "00010101010110001111111111111110";
                        f_reg(164) <= "00010101000101100000000011101011";
                        f_reg(165) <= "10101100000010000000010010000100";
                        f_reg(166) <= "00000001010000010100000000100101";
                        f_reg(167) <= "00000011000011111011000000100101";
                        f_reg(168) <= "00010101010110000000000011100111";
                        f_reg(169) <= "10101100000010100000010010001000";
                        f_reg(170) <= "00000000000010010101010000000011";
                        f_reg(171) <= "00000000000101111100010000000011";
                        f_reg(172) <= "00010101000101100000000011100011";
                        f_reg(173) <= "10101100000010000000010001011000";
                        f_reg(174) <= "00000000110001000011000000100010";
                        f_reg(175) <= "00000010100100101010000000100010";
                        f_reg(176) <= "00100101110010011101010011110111";
                        f_reg(177) <= "00100111100101111101010011110111";
                        f_reg(178) <= "00000000101011010010100000100111";
                        f_reg(179) <= "00000010011110111001100000100111";
                        f_reg(180) <= "00000000000010000010010000000011";
                        f_reg(181) <= "00000000000101101001010000000011";
                        f_reg(182) <= "00101101011011100001011001001101";
                        f_reg(183) <= "00101111001111000001011001001101";
                        f_reg(184) <= "00000001001001110110100000101011";
                        f_reg(185) <= "00000010111101011101100000101011";
                        f_reg(186) <= "00000000010000010101100000100000";
                        f_reg(187) <= "00000010000011111100100000100000";
                        f_reg(188) <= "00000000011000000100100000100100";
                        f_reg(189) <= "00000010001000001011100000100100";
                        f_reg(190) <= "00010101001101110000000011010001";
                        f_reg(191) <= "10101100000010010000010001011100";
                        f_reg(192) <= "00110001100001111000000001111000";
                        f_reg(193) <= "00110011010101011000000001111000";
                        f_reg(194) <= "00000001011011010001000000100011";
                        f_reg(195) <= "00000011001110111000000000100011";
                        f_reg(196) <= "00000001010001000000100000100010";
                        f_reg(197) <= "00000011000100100111100000100010";
                        f_reg(198) <= "00000000110011010001100000101011";
                        f_reg(199) <= "00000010100110111000100000101011";
                        f_reg(200) <= "10001100000010010000010010000000";
                        f_reg(201) <= "10001100000101110000010010000000";
                        f_reg(202) <= "00010101001101111111111111111110";
                        f_reg(203) <= "00000001011010010110000000100101";
                        f_reg(204) <= "00000011001101111101000000100101";
                        f_reg(205) <= "00100101000010101000000100111100";
                        f_reg(206) <= "00100110110110001000000100111100";
                        f_reg(207) <= "00111000101001001100000101001101";
                        f_reg(208) <= "00111010011100101100000101001101";
                        f_reg(209) <= "10001100000010110000010001111100";
                        f_reg(210) <= "10001100000110010000010001111100";
                        f_reg(211) <= "00010101011110011111111111111110";
                        f_reg(212) <= "00010101011110010000000010111011";
                        f_reg(213) <= "10101100000010110000010001100000";
                        f_reg(214) <= "00101100011010010110110111011111";
                        f_reg(215) <= "00101110001101110110110111011111";
                        f_reg(216) <= "00010101100110100000000010110111";
                        f_reg(217) <= "10101100000011000000010001100100";
                        f_reg(218) <= "00010101010110000000000010110101";
                        f_reg(219) <= "10101100000010100000010001101000";
                        f_reg(220) <= "00000001101001000100000000000100";
                        f_reg(221) <= "00000011011100101011000000000100";
                        f_reg(222) <= "00000000111011100010100000101010";
                        f_reg(223) <= "00000010101111001001100000101010";
                        f_reg(224) <= "00000000001010010101100000100110";
                        f_reg(225) <= "00000001111101111100100000100110";
                        f_reg(226) <= "00000000110000110110000000100111";
                        f_reg(227) <= "00000010100100011101000000100111";
                        f_reg(228) <= "00000000000000000000000000000000";
                        f_reg(229) <= "00000000000000000000000000000000";
                        f_reg(230) <= "00010101100110100000000010101001";
                        f_reg(231) <= "10101100000011000000010001101100";
                        f_reg(232) <= "00010100101100110000000010100111";
                        f_reg(233) <= "10101100000001010000010001110000";
                        f_reg(234) <= "00000001000000000101000000100100";
                        f_reg(235) <= "00000010110000001100000000100100";
                        f_reg(236) <= "10001100000001000000010010001000";
                        f_reg(237) <= "10001100000100100000010010001000";
                        f_reg(238) <= "00010100100100101111111111111110";
                        f_reg(239) <= "00000000100000100110100000100010";
                        f_reg(240) <= "00000010010100001101100000100010";
                        f_reg(241) <= "10001100000001110000010010000100";
                        f_reg(242) <= "10001100000101010000010010000100";
                        f_reg(243) <= "00010100111101011111111111111110";
                        f_reg(244) <= "00000000111010110111000000100000";
                        f_reg(245) <= "00000010101110011110000000100000";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00110101010000010111000001000101";
                        f_reg(249) <= "00110111000011110111000001000101";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00000000000000000000000000000000";
                        f_reg(252) <= "00000000001011010100100000101011";
                        f_reg(253) <= "00000001111110111011100000101011";
                        f_reg(254) <= "00010101001101110000000010010001";
                        f_reg(255) <= "10101100000010010000010001110100";
                        f_reg(256) <= "00000000000011100111001111000000";
                        f_reg(257) <= "00000000000111001110001111000000";
                        f_reg(258) <= "00000000000000000000000000000000";
                        f_reg(259) <= "00000000000000000000000000000000";
                        f_reg(260) <= "00010101110111000000000010001011";
                        f_reg(261) <= "10101100000011100000010001111000";
                        f_reg(262) <= "00100011110111011111111100000110";
                        f_reg(263) <= "00010011101000000000000000011101";
                        f_reg(264) <= "00100011110111011111111000001100";
                        f_reg(265) <= "00010011101000000000000000011011";
                        f_reg(266) <= "00100011110111011111110100010010";
                        f_reg(267) <= "00010011101000000000000000011001";
                        f_reg(268) <= "00100011110111101111111111111111";
                        f_reg(269) <= "00100011111111111111111111111111";
                        f_reg(270) <= "00010111110111110000000010000001";
                        f_reg(271) <= "00011111111000001111111101000101";
                        f_reg(272) <= "00010000000000000000000100001100";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "00000000000000000000000000000000";
                        f_reg(287) <= "00000000000000000000000000000000";
                        f_reg(288) <= "00000000000000000000000000000000";
                        f_reg(289) <= "00000000000000000000000000000000";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "10001100000111010000011111100000";
                        f_reg(293) <= "00011111101000000000000000000011";
                        f_reg(294) <= "00100000000111010000000000111100";
                        f_reg(295) <= "00010000000000000000000000000010";
                        f_reg(296) <= "00100000000111010000000000000000";
                        f_reg(297) <= "00010100001011110000000001100110";
                        f_reg(298) <= "10101111101000010000011101101000";
                        f_reg(299) <= "10001100000111010000011111100000";
                        f_reg(300) <= "00011111101000000000000000000011";
                        f_reg(301) <= "00100000000111010000000000111100";
                        f_reg(302) <= "00010000000000000000000000000010";
                        f_reg(303) <= "00100000000111010000000000000000";
                        f_reg(304) <= "00010100010100000000000001011111";
                        f_reg(305) <= "10101111101000100000011101101100";
                        f_reg(306) <= "10001100000111010000011111100000";
                        f_reg(307) <= "00011111101000000000000000000011";
                        f_reg(308) <= "00100000000111010000000000111100";
                        f_reg(309) <= "00010000000000000000000000000010";
                        f_reg(310) <= "00100000000111010000000000000000";
                        f_reg(311) <= "00010100011100010000000001011000";
                        f_reg(312) <= "10101111101000110000011101110000";
                        f_reg(313) <= "10001100000111010000011111100000";
                        f_reg(314) <= "00011111101000000000000000000011";
                        f_reg(315) <= "00100000000111010000000000111100";
                        f_reg(316) <= "00010000000000000000000000000010";
                        f_reg(317) <= "00100000000111010000000000000000";
                        f_reg(318) <= "00010100100100100000000001010001";
                        f_reg(319) <= "10101111101001000000011101110100";
                        f_reg(320) <= "10001100000111010000011111100000";
                        f_reg(321) <= "00011111101000000000000000000011";
                        f_reg(322) <= "00100000000111010000000000111100";
                        f_reg(323) <= "00010000000000000000000000000010";
                        f_reg(324) <= "00100000000111010000000000000000";
                        f_reg(325) <= "00010100101100110000000001001010";
                        f_reg(326) <= "10101111101001010000011101111000";
                        f_reg(327) <= "10001100000111010000011111100000";
                        f_reg(328) <= "00011111101000000000000000000011";
                        f_reg(329) <= "00100000000111010000000000111100";
                        f_reg(330) <= "00010000000000000000000000000010";
                        f_reg(331) <= "00100000000111010000000000000000";
                        f_reg(332) <= "00010100110101000000000001000011";
                        f_reg(333) <= "10101111101001100000011101111100";
                        f_reg(334) <= "10001100000111010000011111100000";
                        f_reg(335) <= "00011111101000000000000000000011";
                        f_reg(336) <= "00100000000111010000000000111100";
                        f_reg(337) <= "00010000000000000000000000000010";
                        f_reg(338) <= "00100000000111010000000000000000";
                        f_reg(339) <= "00010100111101010000000000111100";
                        f_reg(340) <= "10101111101001110000011110000000";
                        f_reg(341) <= "10001100000111010000011111100000";
                        f_reg(342) <= "00011111101000000000000000000011";
                        f_reg(343) <= "00100000000111010000000000111100";
                        f_reg(344) <= "00010000000000000000000000000010";
                        f_reg(345) <= "00100000000111010000000000000000";
                        f_reg(346) <= "00010101000101100000000000110101";
                        f_reg(347) <= "10101111101010000000011110000100";
                        f_reg(348) <= "10001100000111010000011111100000";
                        f_reg(349) <= "00011111101000000000000000000011";
                        f_reg(350) <= "00100000000111010000000000111100";
                        f_reg(351) <= "00010000000000000000000000000010";
                        f_reg(352) <= "00100000000111010000000000000000";
                        f_reg(353) <= "00010101001101110000000000101110";
                        f_reg(354) <= "10101111101010010000011110001000";
                        f_reg(355) <= "10001100000111010000011111100000";
                        f_reg(356) <= "00011111101000000000000000000011";
                        f_reg(357) <= "00100000000111010000000000111100";
                        f_reg(358) <= "00010000000000000000000000000010";
                        f_reg(359) <= "00100000000111010000000000000000";
                        f_reg(360) <= "00010101010110000000000000100111";
                        f_reg(361) <= "10101111101010100000011110001100";
                        f_reg(362) <= "10001100000111010000011111100000";
                        f_reg(363) <= "00011111101000000000000000000011";
                        f_reg(364) <= "00100000000111010000000000111100";
                        f_reg(365) <= "00010000000000000000000000000010";
                        f_reg(366) <= "00100000000111010000000000000000";
                        f_reg(367) <= "00010101011110010000000000100000";
                        f_reg(368) <= "10101111101010110000011110010000";
                        f_reg(369) <= "10001100000111010000011111100000";
                        f_reg(370) <= "00011111101000000000000000000011";
                        f_reg(371) <= "00100000000111010000000000111100";
                        f_reg(372) <= "00010000000000000000000000000010";
                        f_reg(373) <= "00100000000111010000000000000000";
                        f_reg(374) <= "00010101100110100000000000011001";
                        f_reg(375) <= "10101111101011000000011110010100";
                        f_reg(376) <= "10001100000111010000011111100000";
                        f_reg(377) <= "00011111101000000000000000000011";
                        f_reg(378) <= "00100000000111010000000000111100";
                        f_reg(379) <= "00010000000000000000000000000010";
                        f_reg(380) <= "00100000000111010000000000000000";
                        f_reg(381) <= "00010101101110110000000000010010";
                        f_reg(382) <= "10101111101011010000011110011000";
                        f_reg(383) <= "10001100000111010000011111100000";
                        f_reg(384) <= "00011111101000000000000000000011";
                        f_reg(385) <= "00100000000111010000000000111100";
                        f_reg(386) <= "00010000000000000000000000000010";
                        f_reg(387) <= "00100000000111010000000000000000";
                        f_reg(388) <= "00010101110111000000000000001011";
                        f_reg(389) <= "10101111101011100000011110011100";
                        f_reg(390) <= "10001100000111010000011111100000";
                        f_reg(391) <= "00011111101000000000000000000011";
                        f_reg(392) <= "00100000000111010000000000111100";
                        f_reg(393) <= "00010000000000000000000000000010";
                        f_reg(394) <= "00100000000111010000000000000000";
                        f_reg(395) <= "00010111110111110000000000000100";
                        f_reg(396) <= "10101111101111100000011110100000";
                        f_reg(397) <= "10101100000111010000011111100000";
                        f_reg(398) <= "00010000000000001111111101111110";
                        f_reg(399) <= "10001100000111010000011111100000";
                        f_reg(400) <= "10001111101000010000011101101000";
                        f_reg(401) <= "10001100000111010000011111100000";
                        f_reg(402) <= "10001111101011110000011101101000";
                        f_reg(403) <= "00010100001011111111111111111100";
                        f_reg(404) <= "10001100000111010000011111100000";
                        f_reg(405) <= "10001111101000100000011101101100";
                        f_reg(406) <= "10001100000111010000011111100000";
                        f_reg(407) <= "10001111101100000000011101101100";
                        f_reg(408) <= "00010100010100001111111111111100";
                        f_reg(409) <= "10001100000111010000011111100000";
                        f_reg(410) <= "10001111101000110000011101110000";
                        f_reg(411) <= "10001100000111010000011111100000";
                        f_reg(412) <= "10001111101100010000011101110000";
                        f_reg(413) <= "00010100011100011111111111111100";
                        f_reg(414) <= "10001100000111010000011111100000";
                        f_reg(415) <= "10001111101001000000011101110100";
                        f_reg(416) <= "10001100000111010000011111100000";
                        f_reg(417) <= "10001111101100100000011101110100";
                        f_reg(418) <= "00010100100100101111111111111100";
                        f_reg(419) <= "10001100000111010000011111100000";
                        f_reg(420) <= "10001111101001010000011101111000";
                        f_reg(421) <= "10001100000111010000011111100000";
                        f_reg(422) <= "10001111101100110000011101111000";
                        f_reg(423) <= "00010100101100111111111111111100";
                        f_reg(424) <= "10001100000111010000011111100000";
                        f_reg(425) <= "10001111101001100000011101111100";
                        f_reg(426) <= "10001100000111010000011111100000";
                        f_reg(427) <= "10001111101101000000011101111100";
                        f_reg(428) <= "00010100110101001111111111111100";
                        f_reg(429) <= "10001100000111010000011111100000";
                        f_reg(430) <= "10001111101001110000011110000000";
                        f_reg(431) <= "10001100000111010000011111100000";
                        f_reg(432) <= "10001111101101010000011110000000";
                        f_reg(433) <= "00010100111101011111111111111100";
                        f_reg(434) <= "10001100000111010000011111100000";
                        f_reg(435) <= "10001111101010000000011110000100";
                        f_reg(436) <= "10001100000111010000011111100000";
                        f_reg(437) <= "10001111101101100000011110000100";
                        f_reg(438) <= "00010101000101101111111111111100";
                        f_reg(439) <= "10001100000111010000011111100000";
                        f_reg(440) <= "10001111101010010000011110001000";
                        f_reg(441) <= "10001100000111010000011111100000";
                        f_reg(442) <= "10001111101101110000011110001000";
                        f_reg(443) <= "00010101001101111111111111111100";
                        f_reg(444) <= "10001100000111010000011111100000";
                        f_reg(445) <= "10001111101010100000011110001100";
                        f_reg(446) <= "10001100000111010000011111100000";
                        f_reg(447) <= "10001111101110000000011110001100";
                        f_reg(448) <= "00010101010110001111111111111100";
                        f_reg(449) <= "10001100000111010000011111100000";
                        f_reg(450) <= "10001111101010110000011110010000";
                        f_reg(451) <= "10001100000111010000011111100000";
                        f_reg(452) <= "10001111101110010000011110010000";
                        f_reg(453) <= "00010101011110011111111111111100";
                        f_reg(454) <= "10001100000111010000011111100000";
                        f_reg(455) <= "10001111101011000000011110010100";
                        f_reg(456) <= "10001100000111010000011111100000";
                        f_reg(457) <= "10001111101110100000011110010100";
                        f_reg(458) <= "00010101100110101111111111111100";
                        f_reg(459) <= "10001100000111010000011111100000";
                        f_reg(460) <= "10001111101011010000011110011000";
                        f_reg(461) <= "10001100000111010000011111100000";
                        f_reg(462) <= "10001111101110110000011110011000";
                        f_reg(463) <= "00010101101110111111111111111100";
                        f_reg(464) <= "10001100000111010000011111100000";
                        f_reg(465) <= "10001111101011100000011110011100";
                        f_reg(466) <= "10001100000111010000011111100000";
                        f_reg(467) <= "10001111101111000000011110011100";
                        f_reg(468) <= "00010101110111001111111111111100";
                        f_reg(469) <= "10001100000111010000011111100000";
                        f_reg(470) <= "10001111101111100000011110100000";
                        f_reg(471) <= "10001100000111010000011111100000";
                        f_reg(472) <= "10001111101111110000011110100000";
                        f_reg(473) <= "00010111110111111111111111111100";
                        f_reg(474) <= "00010000000000001111111100110010";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000001111100111";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test20_Reg_COMBINED;
