--| LEFT_SHIFT.vhd
--| Implements the left shift function.  Shifts input A by the amount specified by SA.
--|
--| INPUTS:
--| i_A - Data Input
--| i_SA - Shift Amount
--|
--| OUTPUTS:
--| o_Z - Shifted input data (o_Z = i_A << i_SA)
library IEEE;
use IEEE.std_logic_1164.all;

entity LEFT_SHIFT is
	port (i_A	: in  std_logic_vector(31 downto 0);
			i_SA	: in  std_logic_vector(4 downto 0);
			o_Z	: out std_logic_vector(31 downto 0));
end LEFT_SHIFT;

architecture a_LEFT_SHIFT of LEFT_SHIFT is
	-- Declare Components
	component myMUX32_1 is
		port (i_0	: in  std_logic;
				i_1	: in  std_logic;
				i_2	: in  std_logic;
				i_3	: in  std_logic;
				i_4	: in  std_logic;
				i_5	: in  std_logic;
				i_6	: in  std_logic;
				i_7	: in  std_logic;
				i_8	: in  std_logic;
				i_9	: in  std_logic;
				i_10	: in  std_logic;
				i_11	: in  std_logic;
				i_12	: in  std_logic;
				i_13	: in  std_logic;
				i_14	: in  std_logic;
				i_15	: in  std_logic;
				i_16	: in  std_logic;
				i_17	: in  std_logic;
				i_18	: in  std_logic;
				i_19	: in  std_logic;
				i_20	: in  std_logic;
				i_21	: in  std_logic;
				i_22	: in  std_logic;
				i_23	: in  std_logic;
				i_24	: in  std_logic;
				i_25	: in  std_logic;
				i_26	: in  std_logic;
				i_27	: in  std_logic;
				i_28	: in  std_logic;
				i_29	: in  std_logic;
				i_30	: in  std_logic;
				i_31	: in  std_logic;
				i_S	: in  std_logic_vector (4 downto 0);
				o_Z	: out std_logic
				);
	end component;

	-- Declare constants
	constant k_zero : std_logic := '0';

begin	
	u_myMUX_bit31: myMUX32_1
	port map (i_0 => i_A(31),
				 i_1 => i_A(30),
				 i_2 => i_A(29),
				 i_3 => i_A(28),
				 i_4 => i_A(27),
				 i_5 => i_A(26),
				 i_6 => i_A(25),
				 i_7 => i_A(24),
				 i_8 => i_A(23),
				 i_9 => i_A(22),
				 i_10 => i_A(21),
				 i_11 => i_A(20),
				 i_12 => i_A(19),
				 i_13 => i_A(18),
				 i_14 => i_A(17),
				 i_15 => i_A(16),
				 i_16 => i_A(15),
				 i_17 => i_A(14),
				 i_18 => i_A(13),
				 i_19 => i_A(12),
				 i_20 => i_A(11),
				 i_21 => i_A(10),
				 i_22 => i_A(9),
				 i_23 => i_A(8),
				 i_24 => i_A(7),
				 i_25 => i_A(6),
				 i_26 => i_A(5),
				 i_27 => i_A(4),
				 i_28 => i_A(3),
				 i_29 => i_A(2),
				 i_30 => i_A(1),
				 i_31 => i_A(0),
				 i_S => i_SA,
				 o_Z => o_Z(31));
	u_myMUX_bit30: myMUX32_1
	port map (i_0 => i_A(30),
				 i_1 => i_A(29),
				 i_2 => i_A(28),
				 i_3 => i_A(27),
				 i_4 => i_A(26),
				 i_5 => i_A(25),
				 i_6 => i_A(24),
				 i_7 => i_A(23),
				 i_8 => i_A(22),
				 i_9 => i_A(21),
				 i_10 => i_A(20),
				 i_11 => i_A(19),
				 i_12 => i_A(18),
				 i_13 => i_A(17),
				 i_14 => i_A(16),
				 i_15 => i_A(15),
				 i_16 => i_A(14),
				 i_17 => i_A(13),
				 i_18 => i_A(12),
				 i_19 => i_A(11),
				 i_20 => i_A(10),
				 i_21 => i_A(9),
				 i_22 => i_A(8),
				 i_23 => i_A(7),
				 i_24 => i_A(6),
				 i_25 => i_A(5),
				 i_26 => i_A(4),
				 i_27 => i_A(3),
				 i_28 => i_A(2),
				 i_29 => i_A(1),
				 i_30 => i_A(0),
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(30));
				 
	u_myMUX_bit29: myMUX32_1
	port map (i_0 => i_A(29),
				 i_1 => i_A(28),
				 i_2 => i_A(27),
				 i_3 => i_A(26),
				 i_4 => i_A(25),
				 i_5 => i_A(24),
				 i_6 => i_A(23),
				 i_7 => i_A(22),
				 i_8 => i_A(21),
				 i_9 => i_A(20),
				 i_10 => i_A(19),
				 i_11 => i_A(18),
				 i_12 => i_A(17),
				 i_13 => i_A(16),
				 i_14 => i_A(15),
				 i_15 => i_A(14),
				 i_16 => i_A(13),
				 i_17 => i_A(12),
				 i_18 => i_A(11),
				 i_19 => i_A(10),
				 i_20 => i_A(9),
				 i_21 => i_A(8),
				 i_22 => i_A(7),
				 i_23 => i_A(6),
				 i_24 => i_A(5),
				 i_25 => i_A(4),
				 i_26 => i_A(3),
				 i_27 => i_A(2),
				 i_28 => i_A(1),
				 i_29 => i_A(0),
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(29));
	u_myMUX_bit28: myMUX32_1
	port map (i_0 => i_A(28),
				 i_1 => i_A(27),
				 i_2 => i_A(26),
				 i_3 => i_A(25),
				 i_4 => i_A(24),
				 i_5 => i_A(23),
				 i_6 => i_A(22),
				 i_7 => i_A(21),
				 i_8 => i_A(20),
				 i_9 => i_A(19),
				 i_10 => i_A(18),
				 i_11 => i_A(17),
				 i_12 => i_A(16),
				 i_13 => i_A(15),
				 i_14 => i_A(14),
				 i_15 => i_A(13),
				 i_16 => i_A(12),
				 i_17 => i_A(11),
				 i_18 => i_A(10),
				 i_19 => i_A(9),
				 i_20 => i_A(8),
				 i_21 => i_A(7),
				 i_22 => i_A(6),
				 i_23 => i_A(5),
				 i_24 => i_A(4),
				 i_25 => i_A(3),
				 i_26 => i_A(2),
				 i_27 => i_A(1),
				 i_28 => i_A(0),
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(28));
				 
	u_myMUX_bit27: myMUX32_1
	port map (i_0 => i_A(27),
				 i_1 => i_A(26),
				 i_2 => i_A(25),
				 i_3 => i_A(24),
				 i_4 => i_A(23),
				 i_5 => i_A(22),
				 i_6 => i_A(21),
				 i_7 => i_A(20),
				 i_8 => i_A(19),
				 i_9 => i_A(18),
				 i_10 => i_A(17),
				 i_11 => i_A(16),
				 i_12 => i_A(15),
				 i_13 => i_A(14),
				 i_14 => i_A(13),
				 i_15 => i_A(12),
				 i_16 => i_A(11),
				 i_17 => i_A(10),
				 i_18 => i_A(9),
				 i_19 => i_A(8),
				 i_20 => i_A(7),
				 i_21 => i_A(6),
				 i_22 => i_A(5),
				 i_23 => i_A(4),
				 i_24 => i_A(3),
				 i_25 => i_A(2),
				 i_26 => i_A(1),
				 i_27 => i_A(0),
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(27));
	
	u_myMUX_bit26: myMUX32_1
	port map (i_0 => i_A(26),
				 i_1 => i_A(25),
				 i_2 => i_A(24),
				 i_3 => i_A(23),
				 i_4 => i_A(22),
				 i_5 => i_A(21),
				 i_6 => i_A(20),
				 i_7 => i_A(19),
				 i_8 => i_A(18),
				 i_9 => i_A(17),
				 i_10 => i_A(16),
				 i_11 => i_A(15),
				 i_12 => i_A(14),
				 i_13 => i_A(13),
				 i_14 => i_A(12),
				 i_15 => i_A(11),
				 i_16 => i_A(10),
				 i_17 => i_A(9),
				 i_18 => i_A(8),
				 i_19 => i_A(7),
				 i_20 => i_A(6),
				 i_21 => i_A(5),
				 i_22 => i_A(4),
				 i_23 => i_A(3),
				 i_24 => i_A(2),
				 i_25 => i_A(1),
				 i_26 => i_A(0),
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(26));
	
	u_myMUX_bit25: myMUX32_1
	port map (i_0 => i_A(25),
				 i_1 => i_A(24),
				 i_2 => i_A(23),
				 i_3 => i_A(22),
				 i_4 => i_A(21),
				 i_5 => i_A(20),
				 i_6 => i_A(19),
				 i_7 => i_A(18),
				 i_8 => i_A(17),
				 i_9 => i_A(16),
				 i_10 => i_A(15),
				 i_11 => i_A(14),
				 i_12 => i_A(13),
				 i_13 => i_A(12),
				 i_14 => i_A(11),
				 i_15 => i_A(10),
				 i_16 => i_A(9),
				 i_17 => i_A(8),
				 i_18 => i_A(7),
				 i_19 => i_A(6),
				 i_20 => i_A(5),
				 i_21 => i_A(4),
				 i_22 => i_A(3),
				 i_23 => i_A(2),
				 i_24 => i_A(1),
				 i_25 => i_A(0),
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(25));
				 
	u_myMUX_bit24: myMUX32_1
	port map (i_0 => i_A(24),
				 i_1 => i_A(23),
				 i_2 => i_A(22),
				 i_3 => i_A(21),
				 i_4 => i_A(20),
				 i_5 => i_A(19),
				 i_6 => i_A(18),
				 i_7 => i_A(17),
				 i_8 => i_A(16),
				 i_9 => i_A(15),
				 i_10 => i_A(14),
				 i_11 => i_A(13),
				 i_12 => i_A(12),
				 i_13 => i_A(11),
				 i_14 => i_A(10),
				 i_15 => i_A(9),
				 i_16 => i_A(8),
				 i_17 => i_A(7),
				 i_18 => i_A(6),
				 i_19 => i_A(5),
				 i_20 => i_A(4),
				 i_21 => i_A(3),
				 i_22 => i_A(2),
				 i_23 => i_A(1),
				 i_24 => i_A(0),
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(24));
				 
	u_myMUX_bit23: myMUX32_1
	port map (i_0 => i_A(23),
				 i_1 => i_A(22),
				 i_2 => i_A(21),
				 i_3 => i_A(20),
				 i_4 => i_A(19),
				 i_5 => i_A(18),
				 i_6 => i_A(17),
				 i_7 => i_A(16),
				 i_8 => i_A(15),
				 i_9 => i_A(14),
				 i_10 => i_A(13),
				 i_11 => i_A(12),
				 i_12 => i_A(11),
				 i_13 => i_A(10),
				 i_14 => i_A(9),
				 i_15 => i_A(8),
				 i_16 => i_A(7),
				 i_17 => i_A(6),
				 i_18 => i_A(5),
				 i_19 => i_A(4),
				 i_20 => i_A(3),
				 i_21 => i_A(2),
				 i_22 => i_A(1),
				 i_23 => i_A(0),
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(23));
	
	u_myMUX_bit22: myMUX32_1
	port map (i_0 => i_A(22),
				 i_1 => i_A(21),
				 i_2 => i_A(20),
				 i_3 => i_A(19),
				 i_4 => i_A(18),
				 i_5 => i_A(17),
				 i_6 => i_A(16),
				 i_7 => i_A(15),
				 i_8 => i_A(14),
				 i_9 => i_A(13),
				 i_10 => i_A(12),
				 i_11 => i_A(11),
				 i_12 => i_A(10),
				 i_13 => i_A(9),
				 i_14 => i_A(8),
				 i_15 => i_A(7),
				 i_16 => i_A(6),
				 i_17 => i_A(5),
				 i_18 => i_A(4),
				 i_19 => i_A(3),
				 i_20 => i_A(2),
				 i_21 => i_A(1),
				 i_22 => i_A(0),
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(22));
				 
	u_myMUX_bit21: myMUX32_1
	port map (i_0 => i_A(21),
				 i_1 => i_A(20),
				 i_2 => i_A(19),
				 i_3 => i_A(18),
				 i_4 => i_A(17),
				 i_5 => i_A(16),
				 i_6 => i_A(15),
				 i_7 => i_A(14),
				 i_8 => i_A(13),
				 i_9 => i_A(12),
				 i_10 => i_A(11),
				 i_11 => i_A(10),
				 i_12 => i_A(9),
				 i_13 => i_A(8),
				 i_14 => i_A(7),
				 i_15 => i_A(6),
				 i_16 => i_A(5),
				 i_17 => i_A(4),
				 i_18 => i_A(3),
				 i_19 => i_A(2),
				 i_20 => i_A(1),
				 i_21 => i_A(0),
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(21));
				 
	u_myMUX_bit20: myMUX32_1
	port map (i_0 => i_A(20),
				 i_1 => i_A(19),
				 i_2 => i_A(18),
				 i_3 => i_A(17),
				 i_4 => i_A(16),
				 i_5 => i_A(15),
				 i_6 => i_A(14),
				 i_7 => i_A(13),
				 i_8 => i_A(12),
				 i_9 => i_A(11),
				 i_10 => i_A(10),
				 i_11 => i_A(9),
				 i_12 => i_A(8),
				 i_13 => i_A(7),
				 i_14 => i_A(6),
				 i_15 => i_A(5),
				 i_16 => i_A(4),
				 i_17 => i_A(3),
				 i_18 => i_A(2),
				 i_19 => i_A(1),
				 i_20 => i_A(0),
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(20));
				 
	u_myMUX_bit19: myMUX32_1
	port map (i_0 => i_A(19),
				 i_1 => i_A(18),
				 i_2 => i_A(17),
				 i_3 => i_A(16),
				 i_4 => i_A(15),
				 i_5 => i_A(14),
				 i_6 => i_A(13),
				 i_7 => i_A(12),
				 i_8 => i_A(11),
				 i_9 => i_A(10),
				 i_10 => i_A(9),
				 i_11 => i_A(8),
				 i_12 => i_A(7),
				 i_13 => i_A(6),
				 i_14 => i_A(5),
				 i_15 => i_A(4),
				 i_16 => i_A(3),
				 i_17 => i_A(2),
				 i_18 => i_A(1),
				 i_19 => i_A(0),
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(19));
				 
	u_myMUX_bit18: myMUX32_1
	port map (i_0 => i_A(18),
				 i_1 => i_A(17),
				 i_2 => i_A(16),
				 i_3 => i_A(15),
				 i_4 => i_A(14),
				 i_5 => i_A(13),
				 i_6 => i_A(12),
				 i_7 => i_A(11),
				 i_8 => i_A(10),
				 i_9 => i_A(9),
				 i_10 => i_A(8),
				 i_11 => i_A(7),
				 i_12 => i_A(6),
				 i_13 => i_A(5),
				 i_14 => i_A(4),
				 i_15 => i_A(3),
				 i_16 => i_A(2),
				 i_17 => i_A(1),
				 i_18 => i_A(0),
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(18));
				 
	u_myMUX_bit17: myMUX32_1
	port map (i_0 => i_A(17),
				 i_1 => i_A(16),
				 i_2 => i_A(15),
				 i_3 => i_A(14),
				 i_4 => i_A(13),
				 i_5 => i_A(12),
				 i_6 => i_A(11),
				 i_7 => i_A(10),
				 i_8 => i_A(9),
				 i_9 => i_A(8),
				 i_10 => i_A(7),
				 i_11 => i_A(6),
				 i_12 => i_A(5),
				 i_13 => i_A(4),
				 i_14 => i_A(3),
				 i_15 => i_A(2),
				 i_16 => i_A(1),
				 i_17 => i_A(0),
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(17));
				 
	u_myMUX_bit16: myMUX32_1
	port map (i_0 => i_A(16),
				 i_1 => i_A(15),
				 i_2 => i_A(14),
				 i_3 => i_A(13),
				 i_4 => i_A(12),
				 i_5 => i_A(11),
				 i_6 => i_A(10),
				 i_7 => i_A(9),
				 i_8 => i_A(8),
				 i_9 => i_A(7),
				 i_10 => i_A(6),
				 i_11 => i_A(5),
				 i_12 => i_A(4),
				 i_13 => i_A(3),
				 i_14 => i_A(2),
				 i_15 => i_A(1),
				 i_16 => i_A(0),
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(16));
				 
	u_myMUX_bit15: myMUX32_1
	port map (i_0 => i_A(15),
				 i_1 => i_A(14),
				 i_2 => i_A(13),
				 i_3 => i_A(12),
				 i_4 => i_A(11),
				 i_5 => i_A(10),
				 i_6 => i_A(9),
				 i_7 => i_A(8),
				 i_8 => i_A(7),
				 i_9 => i_A(6),
				 i_10 => i_A(5),
				 i_11 => i_A(4),
				 i_12 => i_A(3),
				 i_13 => i_A(2),
				 i_14 => i_A(1),
				 i_15 => i_A(0),
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(15));
				 
	u_myMUX_bit14: myMUX32_1
	port map (i_0 => i_A(14),
				 i_1 => i_A(13),
				 i_2 => i_A(12),
				 i_3 => i_A(11),
				 i_4 => i_A(10),
				 i_5 => i_A(9),
				 i_6 => i_A(8),
				 i_7 => i_A(7),
				 i_8 => i_A(6),
				 i_9 => i_A(5),
				 i_10 => i_A(4),
				 i_11 => i_A(3),
				 i_12 => i_A(2),
				 i_13 => i_A(1),
				 i_14 => i_A(0),
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(14));
				 
	u_myMUX_bit13: myMUX32_1
	port map (i_0 => i_A(13),
				 i_1 => i_A(12),
				 i_2 => i_A(11),
				 i_3 => i_A(10),
				 i_4 => i_A(9),
				 i_5 => i_A(8),
				 i_6 => i_A(7),
				 i_7 => i_A(6),
				 i_8 => i_A(5),
				 i_9 => i_A(4),
				 i_10 => i_A(3),
				 i_11 => i_A(2),
				 i_12 => i_A(1),
				 i_13 => i_A(0),
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(13));
				 
	u_myMUX_bit12: myMUX32_1
	port map (i_0 => i_A(12),
				 i_1 => i_A(11),
				 i_2 => i_A(10),
				 i_3 => i_A(9),
				 i_4 => i_A(8),
				 i_5 => i_A(7),
				 i_6 => i_A(6),
				 i_7 => i_A(5),
				 i_8 => i_A(4),
				 i_9 => i_A(3),
				 i_10 => i_A(2),
				 i_11 => i_A(1),
				 i_12 => i_A(0),
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(12));
				 
	u_myMUX_bit11: myMUX32_1
	port map (i_0 => i_A(11),
				 i_1 => i_A(10),
				 i_2 => i_A(9),
				 i_3 => i_A(8),
				 i_4 => i_A(7),
				 i_5 => i_A(6),
				 i_6 => i_A(5),
				 i_7 => i_A(4),
				 i_8 => i_A(3),
				 i_9 => i_A(2),
				 i_10 => i_A(1),
				 i_11 => i_A(0),
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(11));
				 
	u_myMUX_bit10: myMUX32_1
	port map (i_0 => i_A(10),
				 i_1 => i_A(9),
				 i_2 => i_A(8),
				 i_3 => i_A(7),
				 i_4 => i_A(6),
				 i_5 => i_A(5),
				 i_6 => i_A(4),
				 i_7 => i_A(3),
				 i_8 => i_A(2),
				 i_9 => i_A(1),
				 i_10 => i_A(0),
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(10));
				 
	u_myMUX_bit9: myMUX32_1
	port map (i_0 => i_A(9),
				 i_1 => i_A(8),
				 i_2 => i_A(7),
				 i_3 => i_A(6),
				 i_4 => i_A(5),
				 i_5 => i_A(4),
				 i_6 => i_A(3),
				 i_7 => i_A(2),
				 i_8 => i_A(1),
				 i_9 => i_A(0),
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(9));
				 
	u_myMUX_bit8: myMUX32_1
	port map (i_0 => i_A(8),
				 i_1 => i_A(7),
				 i_2 => i_A(6),
				 i_3 => i_A(5),
				 i_4 => i_A(4),
				 i_5 => i_A(3),
				 i_6 => i_A(2),
				 i_7 => i_A(1),
				 i_8 => i_A(0),
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(8));
				 
	u_myMUX_bit7: myMUX32_1
	port map (i_0 => i_A(7),
				 i_1 => i_A(6),
				 i_2 => i_A(5),
				 i_3 => i_A(4),
				 i_4 => i_A(3),
				 i_5 => i_A(2),
				 i_6 => i_A(1),
				 i_7 => i_A(0),
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(7));
				 
	u_myMUX_bit6: myMUX32_1
	port map (i_0 => i_A(6),
				 i_1 => i_A(5),
				 i_2 => i_A(4),
				 i_3 => i_A(3),
				 i_4 => i_A(2),
				 i_5 => i_A(1),
				 i_6 => i_A(0),
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(6));
				 
	u_myMUX_bit5: myMUX32_1
	port map (i_0 => i_A(5),
				 i_1 => i_A(4),
				 i_2 => i_A(3),
				 i_3 => i_A(2),
				 i_4 => i_A(1),
				 i_5 => i_A(0),
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(5));
				 
	u_myMUX_bit4: myMUX32_1
	port map (i_0 => i_A(4),
				 i_1 => i_A(3),
				 i_2 => i_A(2),
				 i_3 => i_A(1),
				 i_4 => i_A(0),
				 i_5 => k_zero,
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(4));
				 
	u_myMUX_bit3: myMUX32_1
	port map (i_0 => i_A(3),
				 i_1 => i_A(2),
				 i_2 => i_A(1),
				 i_3 => i_A(0),
				 i_4 => k_zero,
				 i_5 => k_zero,
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(3));
				 
	u_myMUX_bit2: myMUX32_1
	port map (i_0 => i_A(2),
				 i_1 => i_A(1),
				 i_2 => i_A(0),
				 i_3 => k_zero,
				 i_4 => k_zero,
				 i_5 => k_zero,
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(2));
				 
	u_myMUX_bit1: myMUX32_1
	port map (i_0 => i_A(1),
				 i_1 => i_A(0),
				 i_2 => k_zero,
				 i_3 => k_zero,
				 i_4 => k_zero,
				 i_5 => k_zero,
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(1));
				 
	u_myMUX_bit0: myMUX32_1
	port map (i_0 => i_A(0),
				 i_1 => k_zero,
				 i_2 => k_zero,
				 i_3 => k_zero,
				 i_4 => k_zero,
				 i_5 => k_zero,
				 i_6 => k_zero,
				 i_7 => k_zero,
				 i_8 => k_zero,
				 i_9 => k_zero,
				 i_10 => k_zero,
				 i_11 => k_zero,
				 i_12 => k_zero,
				 i_13 => k_zero,
				 i_14 => k_zero,
				 i_15 => k_zero,
				 i_16 => k_zero,
				 i_17 => k_zero,
				 i_18 => k_zero,
				 i_19 => k_zero,
				 i_20 => k_zero,
				 i_21 => k_zero,
				 i_22 => k_zero,
				 i_23 => k_zero,
				 i_24 => k_zero,
				 i_25 => k_zero,
				 i_26 => k_zero,
				 i_27 => k_zero,
				 i_28 => k_zero,
				 i_29 => k_zero,
				 i_30 => k_zero,
				 i_31 => k_zero,
				 i_S => i_SA,
				 o_Z => o_Z(0));
end a_LEFT_SHIFT;