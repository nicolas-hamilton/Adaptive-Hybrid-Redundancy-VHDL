--| Test77_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:13:26
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test77_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test77_Reg_COMBINED;

architecture a_Test77_Reg_COMBINED of Test77_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 551) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 551) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100", --  495 - 1980
      "00000000000000000000011111000000", --  496 - 1984
      "00000000000000000000011111000100", --  497 - 1988
      "00000000000000000000011111001000", --  498 - 1992
      "00000000000000000000011111001100", --  499 - 1996
      "00000000000000000000011111010000", --  500 - 2000
      "00000000000000000000011111010100", --  501 - 2004
      "00000000000000000000011111011000", --  502 - 2008
      "00000000000000000000011111011100", --  503 - 2012
      "00000000000000000000011111100000", --  504 - 2016
      "00000000000000000000011111100100", --  505 - 2020
      "00000000000000000000011111101000", --  506 - 2024
      "00000000000000000000011111101100", --  507 - 2028
      "00000000000000000000011111110000", --  508 - 2032
      "00000000000000000000011111110100", --  509 - 2036
      "00000000000000000000011111111000", --  510 - 2040
      "00000000000000000000011111111100", --  511 - 2044
      "00000000000000000000100000000000", --  512 - 2048
      "00000000000000000000100000000100", --  513 - 2052
      "00000000000000000000100000001000", --  514 - 2056
      "00000000000000000000100000001100", --  515 - 2060
      "00000000000000000000100000010000", --  516 - 2064
      "00000000000000000000100000010100", --  517 - 2068
      "00000000000000000000100000011000", --  518 - 2072
      "00000000000000000000100000011100", --  519 - 2076
      "00000000000000000000100000100000", --  520 - 2080
      "00000000000000000000100000100100", --  521 - 2084
      "00000000000000000000100000101000", --  522 - 2088
      "00000000000000000000100000101100", --  523 - 2092
      "00000000000000000000100000110000", --  524 - 2096
      "00000000000000000000100000110100", --  525 - 2100
      "00000000000000000000100000111000", --  526 - 2104
      "00000000000000000000100000111100", --  527 - 2108
      "00000000000000000000100001000000", --  528 - 2112
      "00000000000000000000100001000100", --  529 - 2116
      "00000000000000000000100001001000", --  530 - 2120
      "00000000000000000000100001001100", --  531 - 2124
      "00000000000000000000100001010000", --  532 - 2128
      "00000000000000000000100001010100", --  533 - 2132
      "00000000000000000000100001011000", --  534 - 2136
      "00000000000000000000100001011100", --  535 - 2140
      "00000000000000000000100001100000", --  536 - 2144
      "00000000000000000000100001100100", --  537 - 2148
      "00000000000000000000100001101000", --  538 - 2152
      "00000000000000000000100001101100", --  539 - 2156
      "00000000000000000000100001110000", --  540 - 2160
      "00000000000000000000100001110100", --  541 - 2164
      "00000000000000000000100001111000", --  542 - 2168
      "00000000000000000000100001111100", --  543 - 2172
      "00000000000000000000100010000000", --  544 - 2176
      "00000000000000000000100010000100", --  545 - 2180
      "00000000000000000000100010001000", --  546 - 2184
      "00000000000000000000100010001100", --  547 - 2188
      "00000000000000000000100010010000", --  548 - 2192
      "00000000000000000000100010010100", --  549 - 2196
      "00000000000000000000100010011000");--  550 - 2200

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000011010100100111011", --    2 -    8
      "00000000000000010001000001000000", --    3 -   12
      "00000000001000000001100000100010", --    4 -   16
      "00000000000000000010010101000010", --    5 -   20
      "00000000011000010010100000000100", --    6 -   24
      "00000000011000110011000000100011", --    7 -   28
      "00000000000000010011100000000110", --    8 -   32
      "00101100101010001111110110000111", --    9 -   36
      "00000000111010000100100000100111", --   10 -   40
      "00100000000010100101111010111001", --   11 -   44
      "00000000000000000000000000000000", --   12 -   48
      "00000001001001100101100000100111", --   13 -   52
      "00000001011000010110000000100110", --   14 -   56
      "00000000000000110110100000100111", --   15 -   60
      "00111001000011101111011001100010", --   16 -   64
      "10101100000011100000010010000100", --   17 -   68
      "00110001100011110110000100110011", --   18 -   72
      "00000000010010101000000000100110", --   19 -   76
      "00000001111100001000100000000110", --   20 -   80
      "00000001111000011001000000100110", --   21 -   84
      "00000000000011001001101111000010", --   22 -   88
      "00000000110100000011000000000110", --   23 -   92
      "00000000101010001010000000100101", --   24 -   96
      "00000010010100111010100000000100", --   25 -  100
      "00000001111001011011000000100001", --   26 -  104
      "00000000000001001011100011000011", --   27 -  108
      "00000010100010011100000000100101", --   28 -  112
      "00000010010100011100100000100010", --   29 -  116
      "00000010111101001101000000100011", --   30 -  120
      "00000001101101101101100000100111", --   31 -  124
      "00000000110110111110000000101010", --   32 -  128
      "00000010000011101110100000100101", --   33 -  132
      "00110100110111101101101111000001", --   34 -  136
      "00000011000110000011100000101010", --   35 -  140
      "00000000000000000000000000000000", --   36 -  144
      "00111100000010110110000100010000", --   37 -  148
      "00000000100010110001000000100000", --   38 -  152
      "00000000000000000000000000000000", --   39 -  156
      "00111100000011001110101111111011", --   40 -  160
      "00000000000110000100010010000011", --   41 -  164
      "00000011101101010010100000101010", --   42 -  168
      "00000011100101010100100000100000", --   43 -  172
      "00111001000100011001011011100101", --   44 -  176
      "00000000001011111010000000100001", --   45 -  180
      "00000000000000000000000000000000", --   46 -  184
      "00000000111110100110100000100110", --   47 -  188
      "10101100000001110000010010001000", --   48 -  192
      "00000011001101001011000000100101", --   49 -  196
      "00000011100100011101100000000100", --   50 -  200
      "00000010010010011000000000101011", --   51 -  204
      "00000000000000000000000000000000", --   52 -  208
      "00110000101011101011101000001011", --   53 -  212
      "00000000000011000010001000000000", --   54 -  216
      "00000011011011100101100000100000", --   55 -  220
      "00000010110101101100000000100101", --   56 -  224
      "10101100000100110000010010001100", --   57 -  228
      "00000000000000000000000000000000", --   58 -  232
      "10101100000001100000010010010000", --   59 -  236
      "00000000000110001110100000100010", --   60 -  240
      "00000010111010101010100000100001", --   61 -  244
      "00000000100111010100000000000100", --   62 -  248
      "00000001000111100000100000000100", --   63 -  252
      "00101100010011110000110011111111", --   64 -  256
      "00000000000011011101000110000010", --   65 -  260
      "00000000000000010011100111000010", --   66 -  264
      "00000000011101011100100000101010", --   67 -  268
      "00000000111100001010000000101011", --   68 -  272
      "00000000000110011000111110000011", --   69 -  276
      "00000001111100011110000000100010", --   70 -  280
      "00000000000000000000000000000000", --   71 -  284
      "00101101011100101100001010010100", --   72 -  288
      "10101100000111000000010010010100", --   73 -  292
      "10101100000100100000010010011000", --   74 -  296
      "00000000000000000000000000000000", --   75 -  300
      "00110010100010010100000010101111", --   76 -  304
      "00000000000000000000000000000000", --   77 -  308
      "10101100000110100000010010011100", --   78 -  312
      "10101100000010010000010010100000", --   79 -  316
      "00100011111111111111111111111111", --   80 -  320
      "00011111111000001111111110110001", --   81 -  324
      "00010000000000000000000111010100", --   82 -  328
      "00111100000111100000001111100111", --   83 -  332
      "00111100000111110000001111100111", --   84 -  336
      "00000000000111101111010000000010", --   85 -  340
      "00000000000111111111110000000010", --   86 -  344
      "00111100000000011010100100111011", --   87 -  348
      "00111100000011111010100100111011", --   88 -  352
      "00000000000000010001000001000000", --   89 -  356
      "00000000000011111000000001000000", --   90 -  360
      "00000000001000000001100000100010", --   91 -  364
      "00000001111000001000100000100010", --   92 -  368
      "00000000000000000010010101000010", --   93 -  372
      "00000000000000001001010101000010", --   94 -  376
      "00000000011000010010100000000100", --   95 -  380
      "00000010001011111001100000000100", --   96 -  384
      "00000000011000110011000000100011", --   97 -  388
      "00000010001100011010000000100011", --   98 -  392
      "00000000000000010011100000000110", --   99 -  396
      "00000000000011111010100000000110", --  100 -  400
      "00101100101010001111110110000111", --  101 -  404
      "00101110011101101111110110000111", --  102 -  408
      "00000000111010000100100000100111", --  103 -  412
      "00000010101101101011100000100111", --  104 -  416
      "00100000000010100101111010111001", --  105 -  420
      "00100000000110000101111010111001", --  106 -  424
      "00000000000000000000000000000000", --  107 -  428
      "00000000000000000000000000000000", --  108 -  432
      "00000001001001100101100000100111", --  109 -  436
      "00000010111101001100100000100111", --  110 -  440
      "00000001011000010110000000100110", --  111 -  444
      "00000011001011111101000000100110", --  112 -  448
      "00000000000000110110100000100111", --  113 -  452
      "00000000000100011101100000100111", --  114 -  456
      "00111001000011101111011001100010", --  115 -  460
      "00111010110111001111011001100010", --  116 -  464
      "00010101110111000000000100100100", --  117 -  468
      "10101100000011100000010010000100", --  118 -  472
      "00110001100001110110000100110011", --  119 -  476
      "00110011010101010110000100110011", --  120 -  480
      "00000000010010100101100000100110", --  121 -  484
      "00000010000110001100100000100110", --  122 -  488
      "00000000111010110001000000000110", --  123 -  492
      "00000010101110011000000000000110", --  124 -  496
      "00010100011100010000000100011100", --  125 -  500
      "10101100000000110000010010100100", --  126 -  504
      "00000000111000010001100000100110", --  127 -  508
      "00000010101011111000100000100110", --  128 -  512
      "00010101010110000000000100011000", --  129 -  516
      "10101100000010100000010010101000", --  130 -  520
      "00000000000011000101001111000010", --  131 -  524
      "00000000000110101100001111000010", --  132 -  528
      "00000000110010110011000000000110", --  133 -  532
      "00000010100110011010000000000110", --  134 -  536
      "00000000101010000110000000100101", --  135 -  540
      "00000010011101101101000000100101", --  136 -  544
      "00000000011010100100000000000100", --  137 -  548
      "00000010001110001011000000000100", --  138 -  552
      "00010100110101000000000100001110", --  139 -  556
      "10101100000001100000010010101100", --  140 -  560
      "00000000111001010011000000100001", --  141 -  564
      "00000010101100111010000000100001", --  142 -  568
      "00000000000001000010100011000011", --  143 -  572
      "00000000000100101001100011000011", --  144 -  576
      "00010100101100110000000100001000", --  145 -  580
      "10101100000001010000010010110000", --  146 -  584
      "00000001100010010010100000100101", --  147 -  588
      "00000011010101111001100000100101", --  148 -  592
      "00000000011000100100100000100010", --  149 -  596
      "00000010001100001011100000100010", --  150 -  600
      "10001100000000100000010010110000", --  151 -  604
      "10001100000100000000010010110000", --  152 -  608
      "00010100010100001111111111111110", --  153 -  612
      "00010101010110000000000011111111", --  154 -  616
      "10101100000010100000010010110000", --  155 -  620
      "00000000010011000101000000100011", --  156 -  624
      "00000010000110101100000000100011", --  157 -  628
      "00000001101001100110000000100111", --  158 -  632
      "00000011011101001101000000100111", --  159 -  636
      "10001100000011010000010010101100", --  160 -  640
      "10001100000110110000010010101100", --  161 -  644
      "00010101101110111111111111111110", --  162 -  648
      "00000001101011000011000000101010", --  163 -  652
      "00000011011110101010000000101010", --  164 -  656
      "00000001011011100110000000100101", --  165 -  660
      "00000011001111001101000000100101", --  166 -  664
      "00110101101010111101101111000001", --  167 -  668
      "00110111011110011101101111000001", --  168 -  672
      "00000000101001010111000000101010", --  169 -  676
      "00000010011100111110000000101010", --  170 -  680
      "00000000000000000000000000000000", --  171 -  684
      "00000000000000000000000000000000", --  172 -  688
      "00010101011110010000000011101100", --  173 -  692
      "10101100000010110000010010101100", --  174 -  696
      "00111100000010110110000100010000", --  175 -  700
      "00111100000110010110000100010000", --  176 -  704
      "00010100010100000000000011101000", --  177 -  708
      "10101100000000100000010010110100", --  178 -  712
      "00000000100010110001000000100000", --  179 -  716
      "00000010010110011000000000100000", --  180 -  720
      "00000000000000000000000000000000", --  181 -  724
      "00000000000000000000000000000000", --  182 -  728
      "00111100000001001110101111111011", --  183 -  732
      "00111100000100101110101111111011", --  184 -  736
      "00000000000001010101110010000011", --  185 -  740
      "00000000000100111100110010000011", --  186 -  744
      "00000001100010000010100000101010", --  187 -  748
      "00000011010101101001100000101010", --  188 -  752
      "00000000110010000110000000100000", --  189 -  756
      "00000010100101101101000000100000", --  190 -  760
      "00111001011010001001011011100101", --  191 -  764
      "00111011001101101001011011100101", --  192 -  768
      "00000000001001110101100000100001", --  193 -  772
      "00000001111101011100100000100001", --  194 -  776
      "00000000000000000000000000000000", --  195 -  780
      "00000000000000000000000000000000", --  196 -  784
      "00000001110010100000100000100110", --  197 -  788
      "00000011100110000111100000100110", --  198 -  792
      "00010101110111000000000011010010", --  199 -  796
      "10101100000011100000010010001000", --  200 -  800
      "00000001001010110011100000100101", --  201 -  804
      "00000010111110011010100000100101", --  202 -  808
      "00000000110010000101000000000100", --  203 -  812
      "00000010100101101100000000000100", --  204 -  816
      "00000000011011000111000000101011", --  205 -  820
      "00000010001110101110000000101011", --  206 -  824
      "00000000000000000000000000000000", --  207 -  828
      "00000000000000000000000000000000", --  208 -  832
      "00110000101010011011101000001011", --  209 -  836
      "00110010011101111011101000001011", --  210 -  840
      "00000000000001000101101000000000", --  211 -  844
      "00000000000100101100101000000000", --  212 -  848
      "00000001010010010100000000100000", --  213 -  852
      "00000011000101111011000000100000", --  214 -  856
      "00000000111001110011000000100101", --  215 -  860
      "00000010101101011010000000100101", --  216 -  864
      "10001100000000110000010010110000", --  217 -  868
      "10001100000100010000010010110000", --  218 -  872
      "00010100011100011111111111111110", --  219 -  876
      "00010100011100010000000010111101", --  220 -  880
      "10101100000000110000010010001100", --  221 -  884
      "00000000000000000000000000000000", --  222 -  888
      "00000000000000000000000000000000", --  223 -  892
      "00010101101110110000000010111001", --  224 -  896
      "10101100000011010000010010010000", --  225 -  900
      "00000000000001100110000000100010", --  226 -  904
      "00000000000101001101000000100010", --  227 -  908
      "10001100000001010000010010110100", --  228 -  912
      "10001100000100110000010010110100", --  229 -  916
      "00010100101100111111111111111110", --  230 -  920
      "10001100000001000000010010101000", --  231 -  924
      "10001100000100100000010010101000", --  232 -  928
      "00010100100100101111111111111110", --  233 -  932
      "00000000101001000101000000100001", --  234 -  936
      "00000010011100101100000000100001", --  235 -  940
      "00000001011011000100100000000100", --  236 -  944
      "00000011001110101011100000000100", --  237 -  948
      "10001100000001110000010010101100", --  238 -  952
      "10001100000101010000010010101100", --  239 -  956
      "00010100111101011111111111111110", --  240 -  960
      "00000001001001110001100000000100", --  241 -  964
      "00000010111101011000100000000100", --  242 -  968
      "00101100010011010000110011111111", --  243 -  972
      "00101110000110110000110011111111", --  244 -  976
      "00000000000000010011000110000010", --  245 -  980
      "00000000000011111010000110000010", --  246 -  984
      "00000000000000110010100111000010", --  247 -  988
      "00000000000100011001100111000010", --  248 -  992
      "10001100000001000000010010100100", --  249 -  996
      "10001100000100100000010010100100", --  250 - 1000
      "00010100100100101111111111111110", --  251 - 1004
      "00000000100010100110000000101010", --  252 - 1008
      "00000010010110001101000000101010", --  253 - 1012
      "00000000101011100101100000101011", --  254 - 1016
      "00000010011111001100100000101011", --  255 - 1020
      "00000000000011000011111110000011", --  256 - 1024
      "00000000000110101010111110000011", --  257 - 1028
      "00000001101001110100100000100010", --  258 - 1032
      "00000011011101011011100000100010", --  259 - 1036
      "00000000000000000000000000000000", --  260 - 1040
      "00000000000000000000000000000000", --  261 - 1044
      "00101101000000101100001010010100", --  262 - 1048
      "00101110110100001100001010010100", --  263 - 1052
      "00010101001101110000000010010001", --  264 - 1056
      "10101100000010010000010010010100", --  265 - 1060
      "00010100010100000000000010001111", --  266 - 1064
      "10101100000000100000010010011000", --  267 - 1068
      "00000000000000000000000000000000", --  268 - 1072
      "00000000000000000000000000000000", --  269 - 1076
      "00110001011000010100000010101111", --  270 - 1080
      "00110011001011110100000010101111", --  271 - 1084
      "00000000000000000000000000000000", --  272 - 1088
      "00000000000000000000000000000000", --  273 - 1092
      "00010100110101000000000010000111", --  274 - 1096
      "10101100000001100000010010011100", --  275 - 1100
      "00010100001011110000000010000101", --  276 - 1104
      "10101100000000010000010010100000", --  277 - 1108
      "00100011110111011111111100000110", --  278 - 1112
      "00010011101000000000000000010111", --  279 - 1116
      "00100011110111011111111000001100", --  280 - 1120
      "00010011101000000000000000010101", --  281 - 1124
      "00100011110111011111110100010010", --  282 - 1128
      "00010011101000000000000000010011", --  283 - 1132
      "00100011110111101111111111111111", --  284 - 1136
      "00100011111111111111111111111111", --  285 - 1140
      "00010111110111110000000001111011", --  286 - 1144
      "00011111111000001111111100111000", --  287 - 1148
      "00010000000000000000000100000110", --  288 - 1152
      "00000000000000000000000000000000", --  289 - 1156
      "00000000000000000000000000000000", --  290 - 1160
      "00000000000000000000000000000000", --  291 - 1164
      "00000000000000000000000000000000", --  292 - 1168
      "00000000000000000000000000000000", --  293 - 1172
      "00000000000000000000000000000000", --  294 - 1176
      "00000000000000000000000000000000", --  295 - 1180
      "00000000000000000000000000000000", --  296 - 1184
      "00000000000000000000000000000000", --  297 - 1188
      "00000000000000000000000000000000", --  298 - 1192
      "00000000000000000000000000000000", --  299 - 1196
      "00000000000000000000000000000000", --  300 - 1200
      "00000000000000000000000000000000", --  301 - 1204
      "10001100000111010000100000001100", --  302 - 1208
      "00011111101000000000000000000011", --  303 - 1212
      "00100000000111010000000000111100", --  304 - 1216
      "00010000000000000000000000000010", --  305 - 1220
      "00100000000111010000000000000000", --  306 - 1224
      "00010100001011110000000001100110", --  307 - 1228
      "10101111101000010000011110010100", --  308 - 1232
      "10001100000111010000100000001100", --  309 - 1236
      "00011111101000000000000000000011", --  310 - 1240
      "00100000000111010000000000111100", --  311 - 1244
      "00010000000000000000000000000010", --  312 - 1248
      "00100000000111010000000000000000", --  313 - 1252
      "00010100010100000000000001011111", --  314 - 1256
      "10101111101000100000011110011000", --  315 - 1260
      "10001100000111010000100000001100", --  316 - 1264
      "00011111101000000000000000000011", --  317 - 1268
      "00100000000111010000000000111100", --  318 - 1272
      "00010000000000000000000000000010", --  319 - 1276
      "00100000000111010000000000000000", --  320 - 1280
      "00010100011100010000000001011000", --  321 - 1284
      "10101111101000110000011110011100", --  322 - 1288
      "10001100000111010000100000001100", --  323 - 1292
      "00011111101000000000000000000011", --  324 - 1296
      "00100000000111010000000000111100", --  325 - 1300
      "00010000000000000000000000000010", --  326 - 1304
      "00100000000111010000000000000000", --  327 - 1308
      "00010100100100100000000001010001", --  328 - 1312
      "10101111101001000000011110100000", --  329 - 1316
      "10001100000111010000100000001100", --  330 - 1320
      "00011111101000000000000000000011", --  331 - 1324
      "00100000000111010000000000111100", --  332 - 1328
      "00010000000000000000000000000010", --  333 - 1332
      "00100000000111010000000000000000", --  334 - 1336
      "00010100101100110000000001001010", --  335 - 1340
      "10101111101001010000011110100100", --  336 - 1344
      "10001100000111010000100000001100", --  337 - 1348
      "00011111101000000000000000000011", --  338 - 1352
      "00100000000111010000000000111100", --  339 - 1356
      "00010000000000000000000000000010", --  340 - 1360
      "00100000000111010000000000000000", --  341 - 1364
      "00010100110101000000000001000011", --  342 - 1368
      "10101111101001100000011110101000", --  343 - 1372
      "10001100000111010000100000001100", --  344 - 1376
      "00011111101000000000000000000011", --  345 - 1380
      "00100000000111010000000000111100", --  346 - 1384
      "00010000000000000000000000000010", --  347 - 1388
      "00100000000111010000000000000000", --  348 - 1392
      "00010100111101010000000000111100", --  349 - 1396
      "10101111101001110000011110101100", --  350 - 1400
      "10001100000111010000100000001100", --  351 - 1404
      "00011111101000000000000000000011", --  352 - 1408
      "00100000000111010000000000111100", --  353 - 1412
      "00010000000000000000000000000010", --  354 - 1416
      "00100000000111010000000000000000", --  355 - 1420
      "00010101000101100000000000110101", --  356 - 1424
      "10101111101010000000011110110000", --  357 - 1428
      "10001100000111010000100000001100", --  358 - 1432
      "00011111101000000000000000000011", --  359 - 1436
      "00100000000111010000000000111100", --  360 - 1440
      "00010000000000000000000000000010", --  361 - 1444
      "00100000000111010000000000000000", --  362 - 1448
      "00010101001101110000000000101110", --  363 - 1452
      "10101111101010010000011110110100", --  364 - 1456
      "10001100000111010000100000001100", --  365 - 1460
      "00011111101000000000000000000011", --  366 - 1464
      "00100000000111010000000000111100", --  367 - 1468
      "00010000000000000000000000000010", --  368 - 1472
      "00100000000111010000000000000000", --  369 - 1476
      "00010101010110000000000000100111", --  370 - 1480
      "10101111101010100000011110111000", --  371 - 1484
      "10001100000111010000100000001100", --  372 - 1488
      "00011111101000000000000000000011", --  373 - 1492
      "00100000000111010000000000111100", --  374 - 1496
      "00010000000000000000000000000010", --  375 - 1500
      "00100000000111010000000000000000", --  376 - 1504
      "00010101011110010000000000100000", --  377 - 1508
      "10101111101010110000011110111100", --  378 - 1512
      "10001100000111010000100000001100", --  379 - 1516
      "00011111101000000000000000000011", --  380 - 1520
      "00100000000111010000000000111100", --  381 - 1524
      "00010000000000000000000000000010", --  382 - 1528
      "00100000000111010000000000000000", --  383 - 1532
      "00010101100110100000000000011001", --  384 - 1536
      "10101111101011000000011111000000", --  385 - 1540
      "10001100000111010000100000001100", --  386 - 1544
      "00011111101000000000000000000011", --  387 - 1548
      "00100000000111010000000000111100", --  388 - 1552
      "00010000000000000000000000000010", --  389 - 1556
      "00100000000111010000000000000000", --  390 - 1560
      "00010101101110110000000000010010", --  391 - 1564
      "10101111101011010000011111000100", --  392 - 1568
      "10001100000111010000100000001100", --  393 - 1572
      "00011111101000000000000000000011", --  394 - 1576
      "00100000000111010000000000111100", --  395 - 1580
      "00010000000000000000000000000010", --  396 - 1584
      "00100000000111010000000000000000", --  397 - 1588
      "00010101110111000000000000001011", --  398 - 1592
      "10101111101011100000011111001000", --  399 - 1596
      "10001100000111010000100000001100", --  400 - 1600
      "00011111101000000000000000000011", --  401 - 1604
      "00100000000111010000000000111100", --  402 - 1608
      "00010000000000000000000000000010", --  403 - 1612
      "00100000000111010000000000000000", --  404 - 1616
      "00010111110111110000000000000100", --  405 - 1620
      "10101111101111100000011111001100", --  406 - 1624
      "10101100000111010000100000001100", --  407 - 1628
      "00010000000000001111111110000100", --  408 - 1632
      "10001100000111010000100000001100", --  409 - 1636
      "10001111101000010000011110010100", --  410 - 1640
      "10001100000111010000100000001100", --  411 - 1644
      "10001111101011110000011110010100", --  412 - 1648
      "00010100001011111111111111111100", --  413 - 1652
      "10001100000111010000100000001100", --  414 - 1656
      "10001111101000100000011110011000", --  415 - 1660
      "10001100000111010000100000001100", --  416 - 1664
      "10001111101100000000011110011000", --  417 - 1668
      "00010100010100001111111111111100", --  418 - 1672
      "10001100000111010000100000001100", --  419 - 1676
      "10001111101000110000011110011100", --  420 - 1680
      "10001100000111010000100000001100", --  421 - 1684
      "10001111101100010000011110011100", --  422 - 1688
      "00010100011100011111111111111100", --  423 - 1692
      "10001100000111010000100000001100", --  424 - 1696
      "10001111101001000000011110100000", --  425 - 1700
      "10001100000111010000100000001100", --  426 - 1704
      "10001111101100100000011110100000", --  427 - 1708
      "00010100100100101111111111111100", --  428 - 1712
      "10001100000111010000100000001100", --  429 - 1716
      "10001111101001010000011110100100", --  430 - 1720
      "10001100000111010000100000001100", --  431 - 1724
      "10001111101100110000011110100100", --  432 - 1728
      "00010100101100111111111111111100", --  433 - 1732
      "10001100000111010000100000001100", --  434 - 1736
      "10001111101001100000011110101000", --  435 - 1740
      "10001100000111010000100000001100", --  436 - 1744
      "10001111101101000000011110101000", --  437 - 1748
      "00010100110101001111111111111100", --  438 - 1752
      "10001100000111010000100000001100", --  439 - 1756
      "10001111101001110000011110101100", --  440 - 1760
      "10001100000111010000100000001100", --  441 - 1764
      "10001111101101010000011110101100", --  442 - 1768
      "00010100111101011111111111111100", --  443 - 1772
      "10001100000111010000100000001100", --  444 - 1776
      "10001111101010000000011110110000", --  445 - 1780
      "10001100000111010000100000001100", --  446 - 1784
      "10001111101101100000011110110000", --  447 - 1788
      "00010101000101101111111111111100", --  448 - 1792
      "10001100000111010000100000001100", --  449 - 1796
      "10001111101010010000011110110100", --  450 - 1800
      "10001100000111010000100000001100", --  451 - 1804
      "10001111101101110000011110110100", --  452 - 1808
      "00010101001101111111111111111100", --  453 - 1812
      "10001100000111010000100000001100", --  454 - 1816
      "10001111101010100000011110111000", --  455 - 1820
      "10001100000111010000100000001100", --  456 - 1824
      "10001111101110000000011110111000", --  457 - 1828
      "00010101010110001111111111111100", --  458 - 1832
      "10001100000111010000100000001100", --  459 - 1836
      "10001111101010110000011110111100", --  460 - 1840
      "10001100000111010000100000001100", --  461 - 1844
      "10001111101110010000011110111100", --  462 - 1848
      "00010101011110011111111111111100", --  463 - 1852
      "10001100000111010000100000001100", --  464 - 1856
      "10001111101011000000011111000000", --  465 - 1860
      "10001100000111010000100000001100", --  466 - 1864
      "10001111101110100000011111000000", --  467 - 1868
      "00010101100110101111111111111100", --  468 - 1872
      "10001100000111010000100000001100", --  469 - 1876
      "10001111101011010000011111000100", --  470 - 1880
      "10001100000111010000100000001100", --  471 - 1884
      "10001111101110110000011111000100", --  472 - 1888
      "00010101101110111111111111111100", --  473 - 1892
      "10001100000111010000100000001100", --  474 - 1896
      "10001111101011100000011111001000", --  475 - 1900
      "10001100000111010000100000001100", --  476 - 1904
      "10001111101111000000011111001000", --  477 - 1908
      "00010101110111001111111111111100", --  478 - 1912
      "10001100000111010000100000001100", --  479 - 1916
      "10001111101111100000011111001100", --  480 - 1920
      "10001100000111010000100000001100", --  481 - 1924
      "10001111101111110000011111001100", --  482 - 1928
      "00010111110111111111111111111100", --  483 - 1932
      "00010000000000001111111100111000", --  484 - 1936
      "00000000000000000000000000000000", --  485 - 1940
      "00000000000000000000000000000000", --  486 - 1944
      "00000000000000000000000000000000", --  487 - 1948
      "00000000000000000000000000000000", --  488 - 1952
      "00000000000000000000000000000000", --  489 - 1956
      "00000000000000000000000000000000", --  490 - 1960
      "00000000000000000000000000000000", --  491 - 1964
      "00000000000000000000000000000000", --  492 - 1968
      "00000000000000000000000000000000", --  493 - 1972
      "00000000000000000000000000000000", --  494 - 1976
      "00000000000000000000000000000000", --  495 - 1980
      "00000000000000000000000000000000", --  496 - 1984
      "00000000000000000000000000000000", --  497 - 1988
      "00000000000000000000000000000000", --  498 - 1992
      "00000000000000000000000000000000", --  499 - 1996
      "00000000000000000000000000000000", --  500 - 2000
      "00000000000000000000000000000000", --  501 - 2004
      "00000000000000000000000000000000", --  502 - 2008
      "00000000000000000000000000000000", --  503 - 2012
      "00000000000000000000000000000000", --  504 - 2016
      "00000000000000000000000000000000", --  505 - 2020
      "00000000000000000000000000000000", --  506 - 2024
      "00000000000000000000000000000000", --  507 - 2028
      "00000000000000000000000000000000", --  508 - 2032
      "00000000000000000000000000000000", --  509 - 2036
      "00000000000000000000000000000000", --  510 - 2040
      "00000000000000000000000000000000", --  511 - 2044
      "00000000000000000000000000000000", --  512 - 2048
      "00000000000000000000000000000000", --  513 - 2052
      "00000000000000000000000000000000", --  514 - 2056
      "00000000000000000000001111100111", --  515 - 2060
      "00000000000000000000000000000000", --  516 - 2064
      "00000000000000000000000000000000", --  517 - 2068
      "00000000000000000000000000000000", --  518 - 2072
      "00000000000000000000000000000000", --  519 - 2076
      "00000000000000000000000000000000", --  520 - 2080
      "00000000000000000000000000000000", --  521 - 2084
      "00000000000000000000000000000000", --  522 - 2088
      "00000000000000000000000000000000", --  523 - 2092
      "00000000000000000000000000000000", --  524 - 2096
      "00000000000000000000000000000000", --  525 - 2100
      "00000000000000000000000000000000", --  526 - 2104
      "00000000000000000000000000000000", --  527 - 2108
      "00000000000000000000000000000000", --  528 - 2112
      "00000000000000000000000000000000", --  529 - 2116
      "00000000000000000000000000000000", --  530 - 2120
      "00000000000000000000000000000000", --  531 - 2124
      "00000000000000000000000000000000", --  532 - 2128
      "00000000000000000000000000000000", --  533 - 2132
      "00000000000000000000000000000000", --  534 - 2136
      "00000000000000000000000000000000", --  535 - 2140
      "00000000000000000000000000000000", --  536 - 2144
      "00000000000000000000000000000000", --  537 - 2148
      "00000000000000000000000000000000", --  538 - 2152
      "00000000000000000000000000000000", --  539 - 2156
      "00000000000000000000000000000000", --  540 - 2160
      "00000000000000000000000000000000", --  541 - 2164
      "00000000000000000000000000000000", --  542 - 2168
      "00000000000000000000000000000000", --  543 - 2172
      "00000000000000000000000000000000", --  544 - 2176
      "00000000000000000000000000000000", --  545 - 2180
      "00000000000000000000000000000000", --  546 - 2184
      "00000000000000000000000000000000", --  547 - 2188
      "00000000000000000000000000000000", --  548 - 2192
      "00000000000000000000000000000000", --  549 - 2196
      "00000000000000000000000000000000");--  550 - 2200

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000011010100100111011";
         f_reg(4) <= "00000000000000010001000001000000";
         f_reg(5) <= "00000000001000000001100000100010";
         f_reg(6) <= "00000000000000000010010101000010";
         f_reg(7) <= "00000000011000010010100000000100";
         f_reg(8) <= "00000000011000110011000000100011";
         f_reg(9) <= "00000000000000010011100000000110";
         f_reg(10) <= "00101100101010001111110110000111";
         f_reg(11) <= "00000000111010000100100000100111";
         f_reg(12) <= "00100000000010100101111010111001";
         f_reg(13) <= "00000000000000000000000000000000";
         f_reg(14) <= "00000001001001100101100000100111";
         f_reg(15) <= "00000001011000010110000000100110";
         f_reg(16) <= "00000000000000110110100000100111";
         f_reg(17) <= "00111001000011101111011001100010";
         f_reg(18) <= "10101100000011100000010010000100";
         f_reg(19) <= "00110001100011110110000100110011";
         f_reg(20) <= "00000000010010101000000000100110";
         f_reg(21) <= "00000001111100001000100000000110";
         f_reg(22) <= "00000001111000011001000000100110";
         f_reg(23) <= "00000000000011001001101111000010";
         f_reg(24) <= "00000000110100000011000000000110";
         f_reg(25) <= "00000000101010001010000000100101";
         f_reg(26) <= "00000010010100111010100000000100";
         f_reg(27) <= "00000001111001011011000000100001";
         f_reg(28) <= "00000000000001001011100011000011";
         f_reg(29) <= "00000010100010011100000000100101";
         f_reg(30) <= "00000010010100011100100000100010";
         f_reg(31) <= "00000010111101001101000000100011";
         f_reg(32) <= "00000001101101101101100000100111";
         f_reg(33) <= "00000000110110111110000000101010";
         f_reg(34) <= "00000010000011101110100000100101";
         f_reg(35) <= "00110100110111101101101111000001";
         f_reg(36) <= "00000011000110000011100000101010";
         f_reg(37) <= "00000000000000000000000000000000";
         f_reg(38) <= "00111100000010110110000100010000";
         f_reg(39) <= "00000000100010110001000000100000";
         f_reg(40) <= "00000000000000000000000000000000";
         f_reg(41) <= "00111100000011001110101111111011";
         f_reg(42) <= "00000000000110000100010010000011";
         f_reg(43) <= "00000011101101010010100000101010";
         f_reg(44) <= "00000011100101010100100000100000";
         f_reg(45) <= "00111001000100011001011011100101";
         f_reg(46) <= "00000000001011111010000000100001";
         f_reg(47) <= "00000000000000000000000000000000";
         f_reg(48) <= "00000000111110100110100000100110";
         f_reg(49) <= "10101100000001110000010010001000";
         f_reg(50) <= "00000011001101001011000000100101";
         f_reg(51) <= "00000011100100011101100000000100";
         f_reg(52) <= "00000010010010011000000000101011";
         f_reg(53) <= "00000000000000000000000000000000";
         f_reg(54) <= "00110000101011101011101000001011";
         f_reg(55) <= "00000000000011000010001000000000";
         f_reg(56) <= "00000011011011100101100000100000";
         f_reg(57) <= "00000010110101101100000000100101";
         f_reg(58) <= "10101100000100110000010010001100";
         f_reg(59) <= "00000000000000000000000000000000";
         f_reg(60) <= "10101100000001100000010010010000";
         f_reg(61) <= "00000000000110001110100000100010";
         f_reg(62) <= "00000010111010101010100000100001";
         f_reg(63) <= "00000000100111010100000000000100";
         f_reg(64) <= "00000001000111100000100000000100";
         f_reg(65) <= "00101100010011110000110011111111";
         f_reg(66) <= "00000000000011011101000110000010";
         f_reg(67) <= "00000000000000010011100111000010";
         f_reg(68) <= "00000000011101011100100000101010";
         f_reg(69) <= "00000000111100001010000000101011";
         f_reg(70) <= "00000000000110011000111110000011";
         f_reg(71) <= "00000001111100011110000000100010";
         f_reg(72) <= "00000000000000000000000000000000";
         f_reg(73) <= "00101101011100101100001010010100";
         f_reg(74) <= "10101100000111000000010010010100";
         f_reg(75) <= "10101100000100100000010010011000";
         f_reg(76) <= "00000000000000000000000000000000";
         f_reg(77) <= "00110010100010010100000010101111";
         f_reg(78) <= "00000000000000000000000000000000";
         f_reg(79) <= "10101100000110100000010010011100";
         f_reg(80) <= "10101100000010010000010010100000";
         f_reg(81) <= "00100011111111111111111111111111";
         f_reg(82) <= "00011111111000001111111110110001";
         f_reg(83) <= "00010000000000000000000111010100";
         f_reg(84) <= "00111100000111100000001111100111";
         f_reg(85) <= "00111100000111110000001111100111";
         f_reg(86) <= "00000000000111101111010000000010";
         f_reg(87) <= "00000000000111111111110000000010";
         f_reg(88) <= "00111100000000011010100100111011";
         f_reg(89) <= "00111100000011111010100100111011";
         f_reg(90) <= "00000000000000010001000001000000";
         f_reg(91) <= "00000000000011111000000001000000";
         f_reg(92) <= "00000000001000000001100000100010";
         f_reg(93) <= "00000001111000001000100000100010";
         f_reg(94) <= "00000000000000000010010101000010";
         f_reg(95) <= "00000000000000001001010101000010";
         f_reg(96) <= "00000000011000010010100000000100";
         f_reg(97) <= "00000010001011111001100000000100";
         f_reg(98) <= "00000000011000110011000000100011";
         f_reg(99) <= "00000010001100011010000000100011";
         f_reg(100) <= "00000000000000010011100000000110";
         f_reg(101) <= "00000000000011111010100000000110";
         f_reg(102) <= "00101100101010001111110110000111";
         f_reg(103) <= "00101110011101101111110110000111";
         f_reg(104) <= "00000000111010000100100000100111";
         f_reg(105) <= "00000010101101101011100000100111";
         f_reg(106) <= "00100000000010100101111010111001";
         f_reg(107) <= "00100000000110000101111010111001";
         f_reg(108) <= "00000000000000000000000000000000";
         f_reg(109) <= "00000000000000000000000000000000";
         f_reg(110) <= "00000001001001100101100000100111";
         f_reg(111) <= "00000010111101001100100000100111";
         f_reg(112) <= "00000001011000010110000000100110";
         f_reg(113) <= "00000011001011111101000000100110";
         f_reg(114) <= "00000000000000110110100000100111";
         f_reg(115) <= "00000000000100011101100000100111";
         f_reg(116) <= "00111001000011101111011001100010";
         f_reg(117) <= "00111010110111001111011001100010";
         f_reg(118) <= "00010101110111000000000100100100";
         f_reg(119) <= "10101100000011100000010010000100";
         f_reg(120) <= "00110001100001110110000100110011";
         f_reg(121) <= "00110011010101010110000100110011";
         f_reg(122) <= "00000000010010100101100000100110";
         f_reg(123) <= "00000010000110001100100000100110";
         f_reg(124) <= "00000000111010110001000000000110";
         f_reg(125) <= "00000010101110011000000000000110";
         f_reg(126) <= "00010100011100010000000100011100";
         f_reg(127) <= "10101100000000110000010010100100";
         f_reg(128) <= "00000000111000010001100000100110";
         f_reg(129) <= "00000010101011111000100000100110";
         f_reg(130) <= "00010101010110000000000100011000";
         f_reg(131) <= "10101100000010100000010010101000";
         f_reg(132) <= "00000000000011000101001111000010";
         f_reg(133) <= "00000000000110101100001111000010";
         f_reg(134) <= "00000000110010110011000000000110";
         f_reg(135) <= "00000010100110011010000000000110";
         f_reg(136) <= "00000000101010000110000000100101";
         f_reg(137) <= "00000010011101101101000000100101";
         f_reg(138) <= "00000000011010100100000000000100";
         f_reg(139) <= "00000010001110001011000000000100";
         f_reg(140) <= "00010100110101000000000100001110";
         f_reg(141) <= "10101100000001100000010010101100";
         f_reg(142) <= "00000000111001010011000000100001";
         f_reg(143) <= "00000010101100111010000000100001";
         f_reg(144) <= "00000000000001000010100011000011";
         f_reg(145) <= "00000000000100101001100011000011";
         f_reg(146) <= "00010100101100110000000100001000";
         f_reg(147) <= "10101100000001010000010010110000";
         f_reg(148) <= "00000001100010010010100000100101";
         f_reg(149) <= "00000011010101111001100000100101";
         f_reg(150) <= "00000000011000100100100000100010";
         f_reg(151) <= "00000010001100001011100000100010";
         f_reg(152) <= "10001100000000100000010010110000";
         f_reg(153) <= "10001100000100000000010010110000";
         f_reg(154) <= "00010100010100001111111111111110";
         f_reg(155) <= "00010101010110000000000011111111";
         f_reg(156) <= "10101100000010100000010010110000";
         f_reg(157) <= "00000000010011000101000000100011";
         f_reg(158) <= "00000010000110101100000000100011";
         f_reg(159) <= "00000001101001100110000000100111";
         f_reg(160) <= "00000011011101001101000000100111";
         f_reg(161) <= "10001100000011010000010010101100";
         f_reg(162) <= "10001100000110110000010010101100";
         f_reg(163) <= "00010101101110111111111111111110";
         f_reg(164) <= "00000001101011000011000000101010";
         f_reg(165) <= "00000011011110101010000000101010";
         f_reg(166) <= "00000001011011100110000000100101";
         f_reg(167) <= "00000011001111001101000000100101";
         f_reg(168) <= "00110101101010111101101111000001";
         f_reg(169) <= "00110111011110011101101111000001";
         f_reg(170) <= "00000000101001010111000000101010";
         f_reg(171) <= "00000010011100111110000000101010";
         f_reg(172) <= "00000000000000000000000000000000";
         f_reg(173) <= "00000000000000000000000000000000";
         f_reg(174) <= "00010101011110010000000011101100";
         f_reg(175) <= "10101100000010110000010010101100";
         f_reg(176) <= "00111100000010110110000100010000";
         f_reg(177) <= "00111100000110010110000100010000";
         f_reg(178) <= "00010100010100000000000011101000";
         f_reg(179) <= "10101100000000100000010010110100";
         f_reg(180) <= "00000000100010110001000000100000";
         f_reg(181) <= "00000010010110011000000000100000";
         f_reg(182) <= "00000000000000000000000000000000";
         f_reg(183) <= "00000000000000000000000000000000";
         f_reg(184) <= "00111100000001001110101111111011";
         f_reg(185) <= "00111100000100101110101111111011";
         f_reg(186) <= "00000000000001010101110010000011";
         f_reg(187) <= "00000000000100111100110010000011";
         f_reg(188) <= "00000001100010000010100000101010";
         f_reg(189) <= "00000011010101101001100000101010";
         f_reg(190) <= "00000000110010000110000000100000";
         f_reg(191) <= "00000010100101101101000000100000";
         f_reg(192) <= "00111001011010001001011011100101";
         f_reg(193) <= "00111011001101101001011011100101";
         f_reg(194) <= "00000000001001110101100000100001";
         f_reg(195) <= "00000001111101011100100000100001";
         f_reg(196) <= "00000000000000000000000000000000";
         f_reg(197) <= "00000000000000000000000000000000";
         f_reg(198) <= "00000001110010100000100000100110";
         f_reg(199) <= "00000011100110000111100000100110";
         f_reg(200) <= "00010101110111000000000011010010";
         f_reg(201) <= "10101100000011100000010010001000";
         f_reg(202) <= "00000001001010110011100000100101";
         f_reg(203) <= "00000010111110011010100000100101";
         f_reg(204) <= "00000000110010000101000000000100";
         f_reg(205) <= "00000010100101101100000000000100";
         f_reg(206) <= "00000000011011000111000000101011";
         f_reg(207) <= "00000010001110101110000000101011";
         f_reg(208) <= "00000000000000000000000000000000";
         f_reg(209) <= "00000000000000000000000000000000";
         f_reg(210) <= "00110000101010011011101000001011";
         f_reg(211) <= "00110010011101111011101000001011";
         f_reg(212) <= "00000000000001000101101000000000";
         f_reg(213) <= "00000000000100101100101000000000";
         f_reg(214) <= "00000001010010010100000000100000";
         f_reg(215) <= "00000011000101111011000000100000";
         f_reg(216) <= "00000000111001110011000000100101";
         f_reg(217) <= "00000010101101011010000000100101";
         f_reg(218) <= "10001100000000110000010010110000";
         f_reg(219) <= "10001100000100010000010010110000";
         f_reg(220) <= "00010100011100011111111111111110";
         f_reg(221) <= "00010100011100010000000010111101";
         f_reg(222) <= "10101100000000110000010010001100";
         f_reg(223) <= "00000000000000000000000000000000";
         f_reg(224) <= "00000000000000000000000000000000";
         f_reg(225) <= "00010101101110110000000010111001";
         f_reg(226) <= "10101100000011010000010010010000";
         f_reg(227) <= "00000000000001100110000000100010";
         f_reg(228) <= "00000000000101001101000000100010";
         f_reg(229) <= "10001100000001010000010010110100";
         f_reg(230) <= "10001100000100110000010010110100";
         f_reg(231) <= "00010100101100111111111111111110";
         f_reg(232) <= "10001100000001000000010010101000";
         f_reg(233) <= "10001100000100100000010010101000";
         f_reg(234) <= "00010100100100101111111111111110";
         f_reg(235) <= "00000000101001000101000000100001";
         f_reg(236) <= "00000010011100101100000000100001";
         f_reg(237) <= "00000001011011000100100000000100";
         f_reg(238) <= "00000011001110101011100000000100";
         f_reg(239) <= "10001100000001110000010010101100";
         f_reg(240) <= "10001100000101010000010010101100";
         f_reg(241) <= "00010100111101011111111111111110";
         f_reg(242) <= "00000001001001110001100000000100";
         f_reg(243) <= "00000010111101011000100000000100";
         f_reg(244) <= "00101100010011010000110011111111";
         f_reg(245) <= "00101110000110110000110011111111";
         f_reg(246) <= "00000000000000010011000110000010";
         f_reg(247) <= "00000000000011111010000110000010";
         f_reg(248) <= "00000000000000110010100111000010";
         f_reg(249) <= "00000000000100011001100111000010";
         f_reg(250) <= "10001100000001000000010010100100";
         f_reg(251) <= "10001100000100100000010010100100";
         f_reg(252) <= "00010100100100101111111111111110";
         f_reg(253) <= "00000000100010100110000000101010";
         f_reg(254) <= "00000010010110001101000000101010";
         f_reg(255) <= "00000000101011100101100000101011";
         f_reg(256) <= "00000010011111001100100000101011";
         f_reg(257) <= "00000000000011000011111110000011";
         f_reg(258) <= "00000000000110101010111110000011";
         f_reg(259) <= "00000001101001110100100000100010";
         f_reg(260) <= "00000011011101011011100000100010";
         f_reg(261) <= "00000000000000000000000000000000";
         f_reg(262) <= "00000000000000000000000000000000";
         f_reg(263) <= "00101101000000101100001010010100";
         f_reg(264) <= "00101110110100001100001010010100";
         f_reg(265) <= "00010101001101110000000010010001";
         f_reg(266) <= "10101100000010010000010010010100";
         f_reg(267) <= "00010100010100000000000010001111";
         f_reg(268) <= "10101100000000100000010010011000";
         f_reg(269) <= "00000000000000000000000000000000";
         f_reg(270) <= "00000000000000000000000000000000";
         f_reg(271) <= "00110001011000010100000010101111";
         f_reg(272) <= "00110011001011110100000010101111";
         f_reg(273) <= "00000000000000000000000000000000";
         f_reg(274) <= "00000000000000000000000000000000";
         f_reg(275) <= "00010100110101000000000010000111";
         f_reg(276) <= "10101100000001100000010010011100";
         f_reg(277) <= "00010100001011110000000010000101";
         f_reg(278) <= "10101100000000010000010010100000";
         f_reg(279) <= "00100011110111011111111100000110";
         f_reg(280) <= "00010011101000000000000000010111";
         f_reg(281) <= "00100011110111011111111000001100";
         f_reg(282) <= "00010011101000000000000000010101";
         f_reg(283) <= "00100011110111011111110100010010";
         f_reg(284) <= "00010011101000000000000000010011";
         f_reg(285) <= "00100011110111101111111111111111";
         f_reg(286) <= "00100011111111111111111111111111";
         f_reg(287) <= "00010111110111110000000001111011";
         f_reg(288) <= "00011111111000001111111100111000";
         f_reg(289) <= "00010000000000000000000100000110";
         f_reg(290) <= "00000000000000000000000000000000";
         f_reg(291) <= "00000000000000000000000000000000";
         f_reg(292) <= "00000000000000000000000000000000";
         f_reg(293) <= "00000000000000000000000000000000";
         f_reg(294) <= "00000000000000000000000000000000";
         f_reg(295) <= "00000000000000000000000000000000";
         f_reg(296) <= "00000000000000000000000000000000";
         f_reg(297) <= "00000000000000000000000000000000";
         f_reg(298) <= "00000000000000000000000000000000";
         f_reg(299) <= "00000000000000000000000000000000";
         f_reg(300) <= "00000000000000000000000000000000";
         f_reg(301) <= "00000000000000000000000000000000";
         f_reg(302) <= "00000000000000000000000000000000";
         f_reg(303) <= "10001100000111010000100000001100";
         f_reg(304) <= "00011111101000000000000000000011";
         f_reg(305) <= "00100000000111010000000000111100";
         f_reg(306) <= "00010000000000000000000000000010";
         f_reg(307) <= "00100000000111010000000000000000";
         f_reg(308) <= "00010100001011110000000001100110";
         f_reg(309) <= "10101111101000010000011110010100";
         f_reg(310) <= "10001100000111010000100000001100";
         f_reg(311) <= "00011111101000000000000000000011";
         f_reg(312) <= "00100000000111010000000000111100";
         f_reg(313) <= "00010000000000000000000000000010";
         f_reg(314) <= "00100000000111010000000000000000";
         f_reg(315) <= "00010100010100000000000001011111";
         f_reg(316) <= "10101111101000100000011110011000";
         f_reg(317) <= "10001100000111010000100000001100";
         f_reg(318) <= "00011111101000000000000000000011";
         f_reg(319) <= "00100000000111010000000000111100";
         f_reg(320) <= "00010000000000000000000000000010";
         f_reg(321) <= "00100000000111010000000000000000";
         f_reg(322) <= "00010100011100010000000001011000";
         f_reg(323) <= "10101111101000110000011110011100";
         f_reg(324) <= "10001100000111010000100000001100";
         f_reg(325) <= "00011111101000000000000000000011";
         f_reg(326) <= "00100000000111010000000000111100";
         f_reg(327) <= "00010000000000000000000000000010";
         f_reg(328) <= "00100000000111010000000000000000";
         f_reg(329) <= "00010100100100100000000001010001";
         f_reg(330) <= "10101111101001000000011110100000";
         f_reg(331) <= "10001100000111010000100000001100";
         f_reg(332) <= "00011111101000000000000000000011";
         f_reg(333) <= "00100000000111010000000000111100";
         f_reg(334) <= "00010000000000000000000000000010";
         f_reg(335) <= "00100000000111010000000000000000";
         f_reg(336) <= "00010100101100110000000001001010";
         f_reg(337) <= "10101111101001010000011110100100";
         f_reg(338) <= "10001100000111010000100000001100";
         f_reg(339) <= "00011111101000000000000000000011";
         f_reg(340) <= "00100000000111010000000000111100";
         f_reg(341) <= "00010000000000000000000000000010";
         f_reg(342) <= "00100000000111010000000000000000";
         f_reg(343) <= "00010100110101000000000001000011";
         f_reg(344) <= "10101111101001100000011110101000";
         f_reg(345) <= "10001100000111010000100000001100";
         f_reg(346) <= "00011111101000000000000000000011";
         f_reg(347) <= "00100000000111010000000000111100";
         f_reg(348) <= "00010000000000000000000000000010";
         f_reg(349) <= "00100000000111010000000000000000";
         f_reg(350) <= "00010100111101010000000000111100";
         f_reg(351) <= "10101111101001110000011110101100";
         f_reg(352) <= "10001100000111010000100000001100";
         f_reg(353) <= "00011111101000000000000000000011";
         f_reg(354) <= "00100000000111010000000000111100";
         f_reg(355) <= "00010000000000000000000000000010";
         f_reg(356) <= "00100000000111010000000000000000";
         f_reg(357) <= "00010101000101100000000000110101";
         f_reg(358) <= "10101111101010000000011110110000";
         f_reg(359) <= "10001100000111010000100000001100";
         f_reg(360) <= "00011111101000000000000000000011";
         f_reg(361) <= "00100000000111010000000000111100";
         f_reg(362) <= "00010000000000000000000000000010";
         f_reg(363) <= "00100000000111010000000000000000";
         f_reg(364) <= "00010101001101110000000000101110";
         f_reg(365) <= "10101111101010010000011110110100";
         f_reg(366) <= "10001100000111010000100000001100";
         f_reg(367) <= "00011111101000000000000000000011";
         f_reg(368) <= "00100000000111010000000000111100";
         f_reg(369) <= "00010000000000000000000000000010";
         f_reg(370) <= "00100000000111010000000000000000";
         f_reg(371) <= "00010101010110000000000000100111";
         f_reg(372) <= "10101111101010100000011110111000";
         f_reg(373) <= "10001100000111010000100000001100";
         f_reg(374) <= "00011111101000000000000000000011";
         f_reg(375) <= "00100000000111010000000000111100";
         f_reg(376) <= "00010000000000000000000000000010";
         f_reg(377) <= "00100000000111010000000000000000";
         f_reg(378) <= "00010101011110010000000000100000";
         f_reg(379) <= "10101111101010110000011110111100";
         f_reg(380) <= "10001100000111010000100000001100";
         f_reg(381) <= "00011111101000000000000000000011";
         f_reg(382) <= "00100000000111010000000000111100";
         f_reg(383) <= "00010000000000000000000000000010";
         f_reg(384) <= "00100000000111010000000000000000";
         f_reg(385) <= "00010101100110100000000000011001";
         f_reg(386) <= "10101111101011000000011111000000";
         f_reg(387) <= "10001100000111010000100000001100";
         f_reg(388) <= "00011111101000000000000000000011";
         f_reg(389) <= "00100000000111010000000000111100";
         f_reg(390) <= "00010000000000000000000000000010";
         f_reg(391) <= "00100000000111010000000000000000";
         f_reg(392) <= "00010101101110110000000000010010";
         f_reg(393) <= "10101111101011010000011111000100";
         f_reg(394) <= "10001100000111010000100000001100";
         f_reg(395) <= "00011111101000000000000000000011";
         f_reg(396) <= "00100000000111010000000000111100";
         f_reg(397) <= "00010000000000000000000000000010";
         f_reg(398) <= "00100000000111010000000000000000";
         f_reg(399) <= "00010101110111000000000000001011";
         f_reg(400) <= "10101111101011100000011111001000";
         f_reg(401) <= "10001100000111010000100000001100";
         f_reg(402) <= "00011111101000000000000000000011";
         f_reg(403) <= "00100000000111010000000000111100";
         f_reg(404) <= "00010000000000000000000000000010";
         f_reg(405) <= "00100000000111010000000000000000";
         f_reg(406) <= "00010111110111110000000000000100";
         f_reg(407) <= "10101111101111100000011111001100";
         f_reg(408) <= "10101100000111010000100000001100";
         f_reg(409) <= "00010000000000001111111110000100";
         f_reg(410) <= "10001100000111010000100000001100";
         f_reg(411) <= "10001111101000010000011110010100";
         f_reg(412) <= "10001100000111010000100000001100";
         f_reg(413) <= "10001111101011110000011110010100";
         f_reg(414) <= "00010100001011111111111111111100";
         f_reg(415) <= "10001100000111010000100000001100";
         f_reg(416) <= "10001111101000100000011110011000";
         f_reg(417) <= "10001100000111010000100000001100";
         f_reg(418) <= "10001111101100000000011110011000";
         f_reg(419) <= "00010100010100001111111111111100";
         f_reg(420) <= "10001100000111010000100000001100";
         f_reg(421) <= "10001111101000110000011110011100";
         f_reg(422) <= "10001100000111010000100000001100";
         f_reg(423) <= "10001111101100010000011110011100";
         f_reg(424) <= "00010100011100011111111111111100";
         f_reg(425) <= "10001100000111010000100000001100";
         f_reg(426) <= "10001111101001000000011110100000";
         f_reg(427) <= "10001100000111010000100000001100";
         f_reg(428) <= "10001111101100100000011110100000";
         f_reg(429) <= "00010100100100101111111111111100";
         f_reg(430) <= "10001100000111010000100000001100";
         f_reg(431) <= "10001111101001010000011110100100";
         f_reg(432) <= "10001100000111010000100000001100";
         f_reg(433) <= "10001111101100110000011110100100";
         f_reg(434) <= "00010100101100111111111111111100";
         f_reg(435) <= "10001100000111010000100000001100";
         f_reg(436) <= "10001111101001100000011110101000";
         f_reg(437) <= "10001100000111010000100000001100";
         f_reg(438) <= "10001111101101000000011110101000";
         f_reg(439) <= "00010100110101001111111111111100";
         f_reg(440) <= "10001100000111010000100000001100";
         f_reg(441) <= "10001111101001110000011110101100";
         f_reg(442) <= "10001100000111010000100000001100";
         f_reg(443) <= "10001111101101010000011110101100";
         f_reg(444) <= "00010100111101011111111111111100";
         f_reg(445) <= "10001100000111010000100000001100";
         f_reg(446) <= "10001111101010000000011110110000";
         f_reg(447) <= "10001100000111010000100000001100";
         f_reg(448) <= "10001111101101100000011110110000";
         f_reg(449) <= "00010101000101101111111111111100";
         f_reg(450) <= "10001100000111010000100000001100";
         f_reg(451) <= "10001111101010010000011110110100";
         f_reg(452) <= "10001100000111010000100000001100";
         f_reg(453) <= "10001111101101110000011110110100";
         f_reg(454) <= "00010101001101111111111111111100";
         f_reg(455) <= "10001100000111010000100000001100";
         f_reg(456) <= "10001111101010100000011110111000";
         f_reg(457) <= "10001100000111010000100000001100";
         f_reg(458) <= "10001111101110000000011110111000";
         f_reg(459) <= "00010101010110001111111111111100";
         f_reg(460) <= "10001100000111010000100000001100";
         f_reg(461) <= "10001111101010110000011110111100";
         f_reg(462) <= "10001100000111010000100000001100";
         f_reg(463) <= "10001111101110010000011110111100";
         f_reg(464) <= "00010101011110011111111111111100";
         f_reg(465) <= "10001100000111010000100000001100";
         f_reg(466) <= "10001111101011000000011111000000";
         f_reg(467) <= "10001100000111010000100000001100";
         f_reg(468) <= "10001111101110100000011111000000";
         f_reg(469) <= "00010101100110101111111111111100";
         f_reg(470) <= "10001100000111010000100000001100";
         f_reg(471) <= "10001111101011010000011111000100";
         f_reg(472) <= "10001100000111010000100000001100";
         f_reg(473) <= "10001111101110110000011111000100";
         f_reg(474) <= "00010101101110111111111111111100";
         f_reg(475) <= "10001100000111010000100000001100";
         f_reg(476) <= "10001111101011100000011111001000";
         f_reg(477) <= "10001100000111010000100000001100";
         f_reg(478) <= "10001111101111000000011111001000";
         f_reg(479) <= "00010101110111001111111111111100";
         f_reg(480) <= "10001100000111010000100000001100";
         f_reg(481) <= "10001111101111100000011111001100";
         f_reg(482) <= "10001100000111010000100000001100";
         f_reg(483) <= "10001111101111110000011111001100";
         f_reg(484) <= "00010111110111111111111111111100";
         f_reg(485) <= "00010000000000001111111100111000";
         f_reg(486) <= "00000000000000000000000000000000";
         f_reg(487) <= "00000000000000000000000000000000";
         f_reg(488) <= "00000000000000000000000000000000";
         f_reg(489) <= "00000000000000000000000000000000";
         f_reg(490) <= "00000000000000000000000000000000";
         f_reg(491) <= "00000000000000000000000000000000";
         f_reg(492) <= "00000000000000000000000000000000";
         f_reg(493) <= "00000000000000000000000000000000";
         f_reg(494) <= "00000000000000000000000000000000";
         f_reg(495) <= "00000000000000000000000000000000";
         f_reg(496) <= "00000000000000000000000000000000";
         f_reg(497) <= "00000000000000000000000000000000";
         f_reg(498) <= "00000000000000000000000000000000";
         f_reg(499) <= "00000000000000000000000000000000";
         f_reg(500) <= "00000000000000000000000000000000";
         f_reg(501) <= "00000000000000000000000000000000";
         f_reg(502) <= "00000000000000000000000000000000";
         f_reg(503) <= "00000000000000000000000000000000";
         f_reg(504) <= "00000000000000000000000000000000";
         f_reg(505) <= "00000000000000000000000000000000";
         f_reg(506) <= "00000000000000000000000000000000";
         f_reg(507) <= "00000000000000000000000000000000";
         f_reg(508) <= "00000000000000000000000000000000";
         f_reg(509) <= "00000000000000000000000000000000";
         f_reg(510) <= "00000000000000000000000000000000";
         f_reg(511) <= "00000000000000000000000000000000";
         f_reg(512) <= "00000000000000000000000000000000";
         f_reg(513) <= "00000000000000000000000000000000";
         f_reg(514) <= "00000000000000000000000000000000";
         f_reg(515) <= "00000000000000000000000000000000";
         f_reg(516) <= "00000000000000000000001111100111";
         f_reg(517) <= "00000000000000000000000000000000";
         f_reg(518) <= "00000000000000000000000000000000";
         f_reg(519) <= "00000000000000000000000000000000";
         f_reg(520) <= "00000000000000000000000000000000";
         f_reg(521) <= "00000000000000000000000000000000";
         f_reg(522) <= "00000000000000000000000000000000";
         f_reg(523) <= "00000000000000000000000000000000";
         f_reg(524) <= "00000000000000000000000000000000";
         f_reg(525) <= "00000000000000000000000000000000";
         f_reg(526) <= "00000000000000000000000000000000";
         f_reg(527) <= "00000000000000000000000000000000";
         f_reg(528) <= "00000000000000000000000000000000";
         f_reg(529) <= "00000000000000000000000000000000";
         f_reg(530) <= "00000000000000000000000000000000";
         f_reg(531) <= "00000000000000000000000000000000";
         f_reg(532) <= "00000000000000000000000000000000";
         f_reg(533) <= "00000000000000000000000000000000";
         f_reg(534) <= "00000000000000000000000000000000";
         f_reg(535) <= "00000000000000000000000000000000";
         f_reg(536) <= "00000000000000000000000000000000";
         f_reg(537) <= "00000000000000000000000000000000";
         f_reg(538) <= "00000000000000000000000000000000";
         f_reg(539) <= "00000000000000000000000000000000";
         f_reg(540) <= "00000000000000000000000000000000";
         f_reg(541) <= "00000000000000000000000000000000";
         f_reg(542) <= "00000000000000000000000000000000";
         f_reg(543) <= "00000000000000000000000000000000";
         f_reg(544) <= "00000000000000000000000000000000";
         f_reg(545) <= "00000000000000000000000000000000";
         f_reg(546) <= "00000000000000000000000000000000";
         f_reg(547) <= "00000000000000000000000000000000";
         f_reg(548) <= "00000000000000000000000000000000";
         f_reg(549) <= "00000000000000000000000000000000";
         f_reg(550) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 -22213
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SLL R2 R1 1
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SUB R3 R1 R0
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SRL R4 R0 21
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SLLV R5 R1 R3
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- SUBU R6 R3 R3
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- SRLV R7 R1 R0
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- SLTIU R8 R5 -633
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- NOR R9 R7 R8
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- ADDI R10 R0 24249
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- NOP
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- NOR R11 R9 R6
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- XOR R12 R11 R1
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- NOR R13 R0 R3
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- XORI R14 R8 -2462
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- SW R14 R0 1156
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- ANDI R15 R12 24883
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- XOR R16 R2 R10
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SRLV R17 R16 R15
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- XOR R18 R15 R1
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- SRL R19 R12 15
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- SRLV R6 R16 R6
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- OR R20 R5 R8
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- SLLV R21 R19 R18
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- ADDU R22 R15 R5
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- SRA R23 R4 3
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- OR R24 R20 R9
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- SUB R25 R18 R17
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- SUBU R26 R23 R20
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- NOR R27 R13 R22
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- SLT R28 R6 R27
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- OR R29 R16 R14
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- ORI R30 R6 -9279
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- SLT R7 R24 R24
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- NOP
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- LUI R11 24848
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- ADD R2 R4 R11
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- NOP
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- LUI R12 -5125
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- SRA R8 R24 18
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SLT R5 R29 R21
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- ADD R9 R28 R21
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- XORI R17 R8 -26907
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- ADDU R20 R1 R15
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- NOP
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- XOR R13 R7 R26
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- SW R7 R0 1160
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- OR R22 R25 R20
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SLLV R27 R17 R28
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- SLTU R16 R18 R9
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- NOP
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- ANDI R14 R5 -17909
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SLL R4 R12 8
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- ADD R11 R27 R14
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- OR R24 R22 R22
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- SW R19 R0 1164
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- NOP
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SW R6 R0 1168
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- SUB R29 R0 R24
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- ADDU R21 R23 R10
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- SLLV R8 R29 R4
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- SLLV R1 R30 R8
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- SLTIU R15 R2 3327
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- SRL R26 R13 6
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- SRL R7 R1 7
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- SLT R25 R3 R21
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- SLTU R20 R7 R16
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SRA R17 R25 30
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- SUB R28 R15 R17
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- NOP
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SLTIU R18 R11 -15724
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- SW R28 R0 1172
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- SW R18 R0 1176
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- NOP
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- ANDI R9 R20 16559
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- NOP
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- SW R26 R0 1180
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- SW R9 R0 1184
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- BGTZ R31 -79
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- BEQ R0 R0 468
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- LUI R30 999
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- LUI R31 999
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- LUI R1 -22213
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- LUI R15 -22213
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- SLL R2 R1 1
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- SLL R16 R15 1
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- SUB R3 R1 R0
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- SUB R17 R15 R0
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- SRL R4 R0 21
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- SRL R18 R0 21
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- SLLV R5 R1 R3
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SLLV R19 R15 R17
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SUBU R6 R3 R3
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- SUBU R20 R17 R17
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- SRLV R7 R1 R0
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- SRLV R21 R15 R0
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- SLTIU R8 R5 -633
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SLTIU R22 R19 -633
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- NOR R9 R7 R8
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- NOR R23 R21 R22
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- ADDI R10 R0 24249
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- ADDI R24 R0 24249
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- NOP
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- NOP
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- NOR R11 R9 R6
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- NOR R25 R23 R20
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- XOR R12 R11 R1
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- XOR R26 R25 R15
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- NOR R13 R0 R3
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- NOR R27 R0 R17
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- XORI R14 R8 -2462
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- XORI R28 R22 -2462
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- BNE R14 R28 292
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- SW R14 R0 1156
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- ANDI R7 R12 24883
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- ANDI R21 R26 24883
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- XOR R11 R2 R10
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- XOR R25 R16 R24
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SRLV R2 R11 R7
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- SRLV R16 R25 R21
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- BNE R3 R17 284
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- SW R3 R0 1188
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- XOR R3 R7 R1
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- XOR R17 R21 R15
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- BNE R10 R24 280
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- SW R10 R0 1192
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- SRL R10 R12 15
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- SRL R24 R26 15
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- SRLV R6 R11 R6
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- SRLV R20 R25 R20
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- OR R12 R5 R8
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- OR R26 R19 R22
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SLLV R8 R10 R3
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- SLLV R22 R24 R17
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- BNE R6 R20 270
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- SW R6 R0 1196
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- ADDU R6 R7 R5
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- ADDU R20 R21 R19
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- SRA R5 R4 3
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- SRA R19 R18 3
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- BNE R5 R19 264
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- SW R5 R0 1200
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- OR R5 R12 R9
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- OR R19 R26 R23
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- SUB R9 R3 R2
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- SUB R23 R17 R16
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- LW R2 R0 1200
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- LW R16 R0 1200
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- BNE R2 R16 -2
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- BNE R10 R24 255
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- SW R10 R0 1200
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- SUBU R10 R2 R12
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- SUBU R24 R16 R26
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- NOR R12 R13 R6
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- NOR R26 R27 R20
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- LW R13 R0 1196
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- LW R27 R0 1196
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- BNE R13 R27 -2
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- SLT R6 R13 R12
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- SLT R20 R27 R26
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- OR R12 R11 R14
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- OR R26 R25 R28
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- ORI R11 R13 -9279
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- ORI R25 R27 -9279
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- SLT R14 R5 R5
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- SLT R28 R19 R19
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- NOP
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- NOP
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- BNE R11 R25 236
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- SW R11 R0 1196
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- LUI R11 24848
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- LUI R25 24848
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- BNE R2 R16 232
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- SW R2 R0 1204
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- ADD R2 R4 R11
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- ADD R16 R18 R25
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- NOP
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- NOP
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- LUI R4 -5125
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- LUI R18 -5125
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- SRA R11 R5 18
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- SRA R25 R19 18
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- SLT R5 R12 R8
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- SLT R19 R26 R22
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- ADD R12 R6 R8
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- ADD R26 R20 R22
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- XORI R8 R11 -26907
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- XORI R22 R25 -26907
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- ADDU R11 R1 R7
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- ADDU R25 R15 R21
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- NOP
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- NOP
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- XOR R1 R14 R10
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- XOR R15 R28 R24
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- BNE R14 R28 210
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- SW R14 R0 1160
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- OR R7 R9 R11
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- OR R21 R23 R25
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- SLLV R10 R8 R6
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- SLLV R24 R22 R20
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- SLTU R14 R3 R12
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- SLTU R28 R17 R26
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- NOP
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- NOP
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- ANDI R9 R5 -17909
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- ANDI R23 R19 -17909
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- SLL R11 R4 8
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- SLL R25 R18 8
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- ADD R8 R10 R9
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- ADD R22 R24 R23
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- OR R6 R7 R7
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- OR R20 R21 R21
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- LW R3 R0 1200
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- LW R17 R0 1200
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- BNE R3 R17 -2
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- BNE R3 R17 189
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- SW R3 R0 1164
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- NOP
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- NOP
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- BNE R13 R27 185
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- SW R13 R0 1168
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- SUB R12 R0 R6
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- SUB R26 R0 R20
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- LW R5 R0 1204
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- LW R19 R0 1204
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- BNE R5 R19 -2
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- LW R4 R0 1192
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- LW R18 R0 1192
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- BNE R4 R18 -2
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- ADDU R10 R5 R4
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- ADDU R24 R19 R18
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- SLLV R9 R12 R11
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- SLLV R23 R26 R25
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- LW R7 R0 1196
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- LW R21 R0 1196
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- BNE R7 R21 -2
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- SLLV R3 R7 R9
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- SLLV R17 R21 R23
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- SLTIU R13 R2 3327
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- SLTIU R27 R16 3327
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- SRL R6 R1 6
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- SRL R20 R15 6
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- SRL R5 R3 7
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- SRL R19 R17 7
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- LW R4 R0 1188
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- LW R18 R0 1188
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- BNE R4 R18 -2
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- SLT R12 R4 R10
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- SLT R26 R18 R24
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- SLTU R11 R5 R14
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- SLTU R25 R19 R28
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- SRA R7 R12 30
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- SRA R21 R26 30
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- SUB R9 R13 R7
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- SUB R23 R27 R21
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- NOP
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- NOP
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- SLTIU R2 R8 -15724
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- SLTIU R16 R22 -15724
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- BNE R9 R23 145
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- SW R9 R0 1172
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- BNE R2 R16 143
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- SW R2 R0 1176
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- NOP
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- NOP
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- ANDI R1 R11 16559
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- ANDI R15 R25 16559
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- NOP
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- NOP
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- BNE R6 R20 135
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- SW R6 R0 1180
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- BNE R1 R15 133
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- SW R1 R0 1184
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- BEQ R29 R0 23
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- BEQ R29 R0 21
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- BEQ R29 R0 19
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- BNE R30 R31 123
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- BGTZ R31 -200
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- BEQ R0 R0 262
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- NOP
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- NOP
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- NOP
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- NOP
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- NOP
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- NOP
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- NOP
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- NOP
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- NOP
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- NOP
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- NOP
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- NOP
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- NOP
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- SW R1 R29 1940
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- SW R2 R29 1944
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- SW R3 R29 1948
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- SW R4 R29 1952
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- SW R5 R29 1956
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- SW R6 R29 1960
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- SW R7 R29 1964
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- SW R8 R29 1968
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- SW R9 R29 1972
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- SW R10 R29 1976
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- SW R11 R29 1980
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- SW R12 R29 1984
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- SW R13 R29 1988
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- SW R14 R29 1992
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- SW R30 R29 1996
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- SW R29 R0 2060
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- BEQ R0 R0 -124
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- LW R1 R29 1940
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- LW R15 R29 1940
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- LW R2 R29 1944
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- LW R16 R29 1944
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- LW R3 R29 1948
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- LW R17 R29 1948
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R4 R29 1952
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- LW R18 R29 1952
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- LW R5 R29 1956
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- LW R19 R29 1956
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- LW R6 R29 1960
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- LW R20 R29 1960
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- LW R7 R29 1964
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- LW R21 R29 1964
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- LW R8 R29 1968
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- LW R22 R29 1968
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- LW R9 R29 1972
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- LW R23 R29 1972
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- LW R10 R29 1976
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- LW R24 R29 1976
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- LW R11 R29 1980
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- LW R25 R29 1980
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- LW R12 R29 1984
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- LW R26 R29 1984
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- LW R13 R29 1988
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- LW R27 R29 1988
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- LW R14 R29 1992
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- LW R28 R29 1992
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- LW R30 R29 1996
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- LW R29 R0 2060
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- LW R31 R29 1996
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- BEQ R0 R0 -200
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- NOP
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- NOP
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- NOP
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- NOP
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- NOP
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- NOP
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- NOP
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- NOP
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- NOP
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- NOP
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- NOP
                        f_data <= f_reg(496);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(497) =>
                        -- NOP
                        f_data <= f_reg(497);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(498) =>
                        -- NOP
                        f_data <= f_reg(498);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(499) =>
                        -- NOP
                        f_data <= f_reg(499);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(500) =>
                        -- NOP
                        f_data <= f_reg(500);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(501) =>
                        -- NOP
                        f_data <= f_reg(501);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(502) =>
                        -- NOP
                        f_data <= f_reg(502);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(503) =>
                        -- NOP
                        f_data <= f_reg(503);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(504) =>
                        -- NOP
                        f_data <= f_reg(504);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(505) =>
                        -- NOP
                        f_data <= f_reg(505);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(506) =>
                        -- NOP
                        f_data <= f_reg(506);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(507) =>
                        -- NOP
                        f_data <= f_reg(507);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(508) =>
                        -- NOP
                        f_data <= f_reg(508);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(509) =>
                        -- NOP
                        f_data <= f_reg(509);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(510) =>
                        -- NOP
                        f_data <= f_reg(510);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(511) =>
                        -- NOP
                        f_data <= f_reg(511);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(512) =>
                        -- NOP
                        f_data <= f_reg(512);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(513) =>
                        -- NOP
                        f_data <= f_reg(513);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(514) =>
                        -- NOP
                        f_data <= f_reg(514);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(515) =>
                        -- NOP
                        f_data <= f_reg(515);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(516) =>
                        -- NOP
                        f_data <= f_reg(516);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(517) =>
                        -- NOP
                        f_data <= f_reg(517);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(518) =>
                        -- NOP
                        f_data <= f_reg(518);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(519) =>
                        -- NOP
                        f_data <= f_reg(519);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(520) =>
                        -- NOP
                        f_data <= f_reg(520);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(521) =>
                        -- NOP
                        f_data <= f_reg(521);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(522) =>
                        -- NOP
                        f_data <= f_reg(522);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(523) =>
                        -- NOP
                        f_data <= f_reg(523);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(524) =>
                        -- NOP
                        f_data <= f_reg(524);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(525) =>
                        -- NOP
                        f_data <= f_reg(525);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(526) =>
                        -- NOP
                        f_data <= f_reg(526);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(527) =>
                        -- NOP
                        f_data <= f_reg(527);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(528) =>
                        -- NOP
                        f_data <= f_reg(528);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(529) =>
                        -- NOP
                        f_data <= f_reg(529);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(530) =>
                        -- NOP
                        f_data <= f_reg(530);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(531) =>
                        -- NOP
                        f_data <= f_reg(531);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(532) =>
                        -- NOP
                        f_data <= f_reg(532);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(533) =>
                        -- NOP
                        f_data <= f_reg(533);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(534) =>
                        -- NOP
                        f_data <= f_reg(534);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(535) =>
                        -- NOP
                        f_data <= f_reg(535);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(536) =>
                        -- NOP
                        f_data <= f_reg(536);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(537) =>
                        -- NOP
                        f_data <= f_reg(537);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(538) =>
                        -- NOP
                        f_data <= f_reg(538);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(539) =>
                        -- NOP
                        f_data <= f_reg(539);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(540) =>
                        -- NOP
                        f_data <= f_reg(540);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(541) =>
                        -- NOP
                        f_data <= f_reg(541);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(542) =>
                        -- NOP
                        f_data <= f_reg(542);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(543) =>
                        -- NOP
                        f_data <= f_reg(543);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(544) =>
                        -- NOP
                        f_data <= f_reg(544);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(545) =>
                        -- NOP
                        f_data <= f_reg(545);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(546) =>
                        -- NOP
                        f_data <= f_reg(546);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(547) =>
                        -- NOP
                        f_data <= f_reg(547);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(548) =>
                        -- NOP
                        f_data <= f_reg(548);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(549) =>
                        -- NOP
                        f_data <= f_reg(549);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(550) =>
                        -- NOP
                        f_data <= f_reg(550);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(551) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011010100100111011";
                        f_reg(4) <= "00000000000000010001000001000000";
                        f_reg(5) <= "00000000001000000001100000100010";
                        f_reg(6) <= "00000000000000000010010101000010";
                        f_reg(7) <= "00000000011000010010100000000100";
                        f_reg(8) <= "00000000011000110011000000100011";
                        f_reg(9) <= "00000000000000010011100000000110";
                        f_reg(10) <= "00101100101010001111110110000111";
                        f_reg(11) <= "00000000111010000100100000100111";
                        f_reg(12) <= "00100000000010100101111010111001";
                        f_reg(13) <= "00000000000000000000000000000000";
                        f_reg(14) <= "00000001001001100101100000100111";
                        f_reg(15) <= "00000001011000010110000000100110";
                        f_reg(16) <= "00000000000000110110100000100111";
                        f_reg(17) <= "00111001000011101111011001100010";
                        f_reg(18) <= "10101100000011100000010010000100";
                        f_reg(19) <= "00110001100011110110000100110011";
                        f_reg(20) <= "00000000010010101000000000100110";
                        f_reg(21) <= "00000001111100001000100000000110";
                        f_reg(22) <= "00000001111000011001000000100110";
                        f_reg(23) <= "00000000000011001001101111000010";
                        f_reg(24) <= "00000000110100000011000000000110";
                        f_reg(25) <= "00000000101010001010000000100101";
                        f_reg(26) <= "00000010010100111010100000000100";
                        f_reg(27) <= "00000001111001011011000000100001";
                        f_reg(28) <= "00000000000001001011100011000011";
                        f_reg(29) <= "00000010100010011100000000100101";
                        f_reg(30) <= "00000010010100011100100000100010";
                        f_reg(31) <= "00000010111101001101000000100011";
                        f_reg(32) <= "00000001101101101101100000100111";
                        f_reg(33) <= "00000000110110111110000000101010";
                        f_reg(34) <= "00000010000011101110100000100101";
                        f_reg(35) <= "00110100110111101101101111000001";
                        f_reg(36) <= "00000011000110000011100000101010";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00111100000010110110000100010000";
                        f_reg(39) <= "00000000100010110001000000100000";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "00111100000011001110101111111011";
                        f_reg(42) <= "00000000000110000100010010000011";
                        f_reg(43) <= "00000011101101010010100000101010";
                        f_reg(44) <= "00000011100101010100100000100000";
                        f_reg(45) <= "00111001000100011001011011100101";
                        f_reg(46) <= "00000000001011111010000000100001";
                        f_reg(47) <= "00000000000000000000000000000000";
                        f_reg(48) <= "00000000111110100110100000100110";
                        f_reg(49) <= "10101100000001110000010010001000";
                        f_reg(50) <= "00000011001101001011000000100101";
                        f_reg(51) <= "00000011100100011101100000000100";
                        f_reg(52) <= "00000010010010011000000000101011";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00110000101011101011101000001011";
                        f_reg(55) <= "00000000000011000010001000000000";
                        f_reg(56) <= "00000011011011100101100000100000";
                        f_reg(57) <= "00000010110101101100000000100101";
                        f_reg(58) <= "10101100000100110000010010001100";
                        f_reg(59) <= "00000000000000000000000000000000";
                        f_reg(60) <= "10101100000001100000010010010000";
                        f_reg(61) <= "00000000000110001110100000100010";
                        f_reg(62) <= "00000010111010101010100000100001";
                        f_reg(63) <= "00000000100111010100000000000100";
                        f_reg(64) <= "00000001000111100000100000000100";
                        f_reg(65) <= "00101100010011110000110011111111";
                        f_reg(66) <= "00000000000011011101000110000010";
                        f_reg(67) <= "00000000000000010011100111000010";
                        f_reg(68) <= "00000000011101011100100000101010";
                        f_reg(69) <= "00000000111100001010000000101011";
                        f_reg(70) <= "00000000000110011000111110000011";
                        f_reg(71) <= "00000001111100011110000000100010";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "00101101011100101100001010010100";
                        f_reg(74) <= "10101100000111000000010010010100";
                        f_reg(75) <= "10101100000100100000010010011000";
                        f_reg(76) <= "00000000000000000000000000000000";
                        f_reg(77) <= "00110010100010010100000010101111";
                        f_reg(78) <= "00000000000000000000000000000000";
                        f_reg(79) <= "10101100000110100000010010011100";
                        f_reg(80) <= "10101100000010010000010010100000";
                        f_reg(81) <= "00100011111111111111111111111111";
                        f_reg(82) <= "00011111111000001111111110110001";
                        f_reg(83) <= "00010000000000000000000111010100";
                        f_reg(84) <= "00111100000111100000001111100111";
                        f_reg(85) <= "00111100000111110000001111100111";
                        f_reg(86) <= "00000000000111101111010000000010";
                        f_reg(87) <= "00000000000111111111110000000010";
                        f_reg(88) <= "00111100000000011010100100111011";
                        f_reg(89) <= "00111100000011111010100100111011";
                        f_reg(90) <= "00000000000000010001000001000000";
                        f_reg(91) <= "00000000000011111000000001000000";
                        f_reg(92) <= "00000000001000000001100000100010";
                        f_reg(93) <= "00000001111000001000100000100010";
                        f_reg(94) <= "00000000000000000010010101000010";
                        f_reg(95) <= "00000000000000001001010101000010";
                        f_reg(96) <= "00000000011000010010100000000100";
                        f_reg(97) <= "00000010001011111001100000000100";
                        f_reg(98) <= "00000000011000110011000000100011";
                        f_reg(99) <= "00000010001100011010000000100011";
                        f_reg(100) <= "00000000000000010011100000000110";
                        f_reg(101) <= "00000000000011111010100000000110";
                        f_reg(102) <= "00101100101010001111110110000111";
                        f_reg(103) <= "00101110011101101111110110000111";
                        f_reg(104) <= "00000000111010000100100000100111";
                        f_reg(105) <= "00000010101101101011100000100111";
                        f_reg(106) <= "00100000000010100101111010111001";
                        f_reg(107) <= "00100000000110000101111010111001";
                        f_reg(108) <= "00000000000000000000000000000000";
                        f_reg(109) <= "00000000000000000000000000000000";
                        f_reg(110) <= "00000001001001100101100000100111";
                        f_reg(111) <= "00000010111101001100100000100111";
                        f_reg(112) <= "00000001011000010110000000100110";
                        f_reg(113) <= "00000011001011111101000000100110";
                        f_reg(114) <= "00000000000000110110100000100111";
                        f_reg(115) <= "00000000000100011101100000100111";
                        f_reg(116) <= "00111001000011101111011001100010";
                        f_reg(117) <= "00111010110111001111011001100010";
                        f_reg(118) <= "00010101110111000000000100100100";
                        f_reg(119) <= "10101100000011100000010010000100";
                        f_reg(120) <= "00110001100001110110000100110011";
                        f_reg(121) <= "00110011010101010110000100110011";
                        f_reg(122) <= "00000000010010100101100000100110";
                        f_reg(123) <= "00000010000110001100100000100110";
                        f_reg(124) <= "00000000111010110001000000000110";
                        f_reg(125) <= "00000010101110011000000000000110";
                        f_reg(126) <= "00010100011100010000000100011100";
                        f_reg(127) <= "10101100000000110000010010100100";
                        f_reg(128) <= "00000000111000010001100000100110";
                        f_reg(129) <= "00000010101011111000100000100110";
                        f_reg(130) <= "00010101010110000000000100011000";
                        f_reg(131) <= "10101100000010100000010010101000";
                        f_reg(132) <= "00000000000011000101001111000010";
                        f_reg(133) <= "00000000000110101100001111000010";
                        f_reg(134) <= "00000000110010110011000000000110";
                        f_reg(135) <= "00000010100110011010000000000110";
                        f_reg(136) <= "00000000101010000110000000100101";
                        f_reg(137) <= "00000010011101101101000000100101";
                        f_reg(138) <= "00000000011010100100000000000100";
                        f_reg(139) <= "00000010001110001011000000000100";
                        f_reg(140) <= "00010100110101000000000100001110";
                        f_reg(141) <= "10101100000001100000010010101100";
                        f_reg(142) <= "00000000111001010011000000100001";
                        f_reg(143) <= "00000010101100111010000000100001";
                        f_reg(144) <= "00000000000001000010100011000011";
                        f_reg(145) <= "00000000000100101001100011000011";
                        f_reg(146) <= "00010100101100110000000100001000";
                        f_reg(147) <= "10101100000001010000010010110000";
                        f_reg(148) <= "00000001100010010010100000100101";
                        f_reg(149) <= "00000011010101111001100000100101";
                        f_reg(150) <= "00000000011000100100100000100010";
                        f_reg(151) <= "00000010001100001011100000100010";
                        f_reg(152) <= "10001100000000100000010010110000";
                        f_reg(153) <= "10001100000100000000010010110000";
                        f_reg(154) <= "00010100010100001111111111111110";
                        f_reg(155) <= "00010101010110000000000011111111";
                        f_reg(156) <= "10101100000010100000010010110000";
                        f_reg(157) <= "00000000010011000101000000100011";
                        f_reg(158) <= "00000010000110101100000000100011";
                        f_reg(159) <= "00000001101001100110000000100111";
                        f_reg(160) <= "00000011011101001101000000100111";
                        f_reg(161) <= "10001100000011010000010010101100";
                        f_reg(162) <= "10001100000110110000010010101100";
                        f_reg(163) <= "00010101101110111111111111111110";
                        f_reg(164) <= "00000001101011000011000000101010";
                        f_reg(165) <= "00000011011110101010000000101010";
                        f_reg(166) <= "00000001011011100110000000100101";
                        f_reg(167) <= "00000011001111001101000000100101";
                        f_reg(168) <= "00110101101010111101101111000001";
                        f_reg(169) <= "00110111011110011101101111000001";
                        f_reg(170) <= "00000000101001010111000000101010";
                        f_reg(171) <= "00000010011100111110000000101010";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00000000000000000000000000000000";
                        f_reg(174) <= "00010101011110010000000011101100";
                        f_reg(175) <= "10101100000010110000010010101100";
                        f_reg(176) <= "00111100000010110110000100010000";
                        f_reg(177) <= "00111100000110010110000100010000";
                        f_reg(178) <= "00010100010100000000000011101000";
                        f_reg(179) <= "10101100000000100000010010110100";
                        f_reg(180) <= "00000000100010110001000000100000";
                        f_reg(181) <= "00000010010110011000000000100000";
                        f_reg(182) <= "00000000000000000000000000000000";
                        f_reg(183) <= "00000000000000000000000000000000";
                        f_reg(184) <= "00111100000001001110101111111011";
                        f_reg(185) <= "00111100000100101110101111111011";
                        f_reg(186) <= "00000000000001010101110010000011";
                        f_reg(187) <= "00000000000100111100110010000011";
                        f_reg(188) <= "00000001100010000010100000101010";
                        f_reg(189) <= "00000011010101101001100000101010";
                        f_reg(190) <= "00000000110010000110000000100000";
                        f_reg(191) <= "00000010100101101101000000100000";
                        f_reg(192) <= "00111001011010001001011011100101";
                        f_reg(193) <= "00111011001101101001011011100101";
                        f_reg(194) <= "00000000001001110101100000100001";
                        f_reg(195) <= "00000001111101011100100000100001";
                        f_reg(196) <= "00000000000000000000000000000000";
                        f_reg(197) <= "00000000000000000000000000000000";
                        f_reg(198) <= "00000001110010100000100000100110";
                        f_reg(199) <= "00000011100110000111100000100110";
                        f_reg(200) <= "00010101110111000000000011010010";
                        f_reg(201) <= "10101100000011100000010010001000";
                        f_reg(202) <= "00000001001010110011100000100101";
                        f_reg(203) <= "00000010111110011010100000100101";
                        f_reg(204) <= "00000000110010000101000000000100";
                        f_reg(205) <= "00000010100101101100000000000100";
                        f_reg(206) <= "00000000011011000111000000101011";
                        f_reg(207) <= "00000010001110101110000000101011";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00110000101010011011101000001011";
                        f_reg(211) <= "00110010011101111011101000001011";
                        f_reg(212) <= "00000000000001000101101000000000";
                        f_reg(213) <= "00000000000100101100101000000000";
                        f_reg(214) <= "00000001010010010100000000100000";
                        f_reg(215) <= "00000011000101111011000000100000";
                        f_reg(216) <= "00000000111001110011000000100101";
                        f_reg(217) <= "00000010101101011010000000100101";
                        f_reg(218) <= "10001100000000110000010010110000";
                        f_reg(219) <= "10001100000100010000010010110000";
                        f_reg(220) <= "00010100011100011111111111111110";
                        f_reg(221) <= "00010100011100010000000010111101";
                        f_reg(222) <= "10101100000000110000010010001100";
                        f_reg(223) <= "00000000000000000000000000000000";
                        f_reg(224) <= "00000000000000000000000000000000";
                        f_reg(225) <= "00010101101110110000000010111001";
                        f_reg(226) <= "10101100000011010000010010010000";
                        f_reg(227) <= "00000000000001100110000000100010";
                        f_reg(228) <= "00000000000101001101000000100010";
                        f_reg(229) <= "10001100000001010000010010110100";
                        f_reg(230) <= "10001100000100110000010010110100";
                        f_reg(231) <= "00010100101100111111111111111110";
                        f_reg(232) <= "10001100000001000000010010101000";
                        f_reg(233) <= "10001100000100100000010010101000";
                        f_reg(234) <= "00010100100100101111111111111110";
                        f_reg(235) <= "00000000101001000101000000100001";
                        f_reg(236) <= "00000010011100101100000000100001";
                        f_reg(237) <= "00000001011011000100100000000100";
                        f_reg(238) <= "00000011001110101011100000000100";
                        f_reg(239) <= "10001100000001110000010010101100";
                        f_reg(240) <= "10001100000101010000010010101100";
                        f_reg(241) <= "00010100111101011111111111111110";
                        f_reg(242) <= "00000001001001110001100000000100";
                        f_reg(243) <= "00000010111101011000100000000100";
                        f_reg(244) <= "00101100010011010000110011111111";
                        f_reg(245) <= "00101110000110110000110011111111";
                        f_reg(246) <= "00000000000000010011000110000010";
                        f_reg(247) <= "00000000000011111010000110000010";
                        f_reg(248) <= "00000000000000110010100111000010";
                        f_reg(249) <= "00000000000100011001100111000010";
                        f_reg(250) <= "10001100000001000000010010100100";
                        f_reg(251) <= "10001100000100100000010010100100";
                        f_reg(252) <= "00010100100100101111111111111110";
                        f_reg(253) <= "00000000100010100110000000101010";
                        f_reg(254) <= "00000010010110001101000000101010";
                        f_reg(255) <= "00000000101011100101100000101011";
                        f_reg(256) <= "00000010011111001100100000101011";
                        f_reg(257) <= "00000000000011000011111110000011";
                        f_reg(258) <= "00000000000110101010111110000011";
                        f_reg(259) <= "00000001101001110100100000100010";
                        f_reg(260) <= "00000011011101011011100000100010";
                        f_reg(261) <= "00000000000000000000000000000000";
                        f_reg(262) <= "00000000000000000000000000000000";
                        f_reg(263) <= "00101101000000101100001010010100";
                        f_reg(264) <= "00101110110100001100001010010100";
                        f_reg(265) <= "00010101001101110000000010010001";
                        f_reg(266) <= "10101100000010010000010010010100";
                        f_reg(267) <= "00010100010100000000000010001111";
                        f_reg(268) <= "10101100000000100000010010011000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00110001011000010100000010101111";
                        f_reg(272) <= "00110011001011110100000010101111";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00010100110101000000000010000111";
                        f_reg(276) <= "10101100000001100000010010011100";
                        f_reg(277) <= "00010100001011110000000010000101";
                        f_reg(278) <= "10101100000000010000010010100000";
                        f_reg(279) <= "00100011110111011111111100000110";
                        f_reg(280) <= "00010011101000000000000000010111";
                        f_reg(281) <= "00100011110111011111111000001100";
                        f_reg(282) <= "00010011101000000000000000010101";
                        f_reg(283) <= "00100011110111011111110100010010";
                        f_reg(284) <= "00010011101000000000000000010011";
                        f_reg(285) <= "00100011110111101111111111111111";
                        f_reg(286) <= "00100011111111111111111111111111";
                        f_reg(287) <= "00010111110111110000000001111011";
                        f_reg(288) <= "00011111111000001111111100111000";
                        f_reg(289) <= "00010000000000000000000100000110";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "00000000000000000000000000000000";
                        f_reg(293) <= "00000000000000000000000000000000";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "10001100000111010000100000001100";
                        f_reg(304) <= "00011111101000000000000000000011";
                        f_reg(305) <= "00100000000111010000000000111100";
                        f_reg(306) <= "00010000000000000000000000000010";
                        f_reg(307) <= "00100000000111010000000000000000";
                        f_reg(308) <= "00010100001011110000000001100110";
                        f_reg(309) <= "10101111101000010000011110010100";
                        f_reg(310) <= "10001100000111010000100000001100";
                        f_reg(311) <= "00011111101000000000000000000011";
                        f_reg(312) <= "00100000000111010000000000111100";
                        f_reg(313) <= "00010000000000000000000000000010";
                        f_reg(314) <= "00100000000111010000000000000000";
                        f_reg(315) <= "00010100010100000000000001011111";
                        f_reg(316) <= "10101111101000100000011110011000";
                        f_reg(317) <= "10001100000111010000100000001100";
                        f_reg(318) <= "00011111101000000000000000000011";
                        f_reg(319) <= "00100000000111010000000000111100";
                        f_reg(320) <= "00010000000000000000000000000010";
                        f_reg(321) <= "00100000000111010000000000000000";
                        f_reg(322) <= "00010100011100010000000001011000";
                        f_reg(323) <= "10101111101000110000011110011100";
                        f_reg(324) <= "10001100000111010000100000001100";
                        f_reg(325) <= "00011111101000000000000000000011";
                        f_reg(326) <= "00100000000111010000000000111100";
                        f_reg(327) <= "00010000000000000000000000000010";
                        f_reg(328) <= "00100000000111010000000000000000";
                        f_reg(329) <= "00010100100100100000000001010001";
                        f_reg(330) <= "10101111101001000000011110100000";
                        f_reg(331) <= "10001100000111010000100000001100";
                        f_reg(332) <= "00011111101000000000000000000011";
                        f_reg(333) <= "00100000000111010000000000111100";
                        f_reg(334) <= "00010000000000000000000000000010";
                        f_reg(335) <= "00100000000111010000000000000000";
                        f_reg(336) <= "00010100101100110000000001001010";
                        f_reg(337) <= "10101111101001010000011110100100";
                        f_reg(338) <= "10001100000111010000100000001100";
                        f_reg(339) <= "00011111101000000000000000000011";
                        f_reg(340) <= "00100000000111010000000000111100";
                        f_reg(341) <= "00010000000000000000000000000010";
                        f_reg(342) <= "00100000000111010000000000000000";
                        f_reg(343) <= "00010100110101000000000001000011";
                        f_reg(344) <= "10101111101001100000011110101000";
                        f_reg(345) <= "10001100000111010000100000001100";
                        f_reg(346) <= "00011111101000000000000000000011";
                        f_reg(347) <= "00100000000111010000000000111100";
                        f_reg(348) <= "00010000000000000000000000000010";
                        f_reg(349) <= "00100000000111010000000000000000";
                        f_reg(350) <= "00010100111101010000000000111100";
                        f_reg(351) <= "10101111101001110000011110101100";
                        f_reg(352) <= "10001100000111010000100000001100";
                        f_reg(353) <= "00011111101000000000000000000011";
                        f_reg(354) <= "00100000000111010000000000111100";
                        f_reg(355) <= "00010000000000000000000000000010";
                        f_reg(356) <= "00100000000111010000000000000000";
                        f_reg(357) <= "00010101000101100000000000110101";
                        f_reg(358) <= "10101111101010000000011110110000";
                        f_reg(359) <= "10001100000111010000100000001100";
                        f_reg(360) <= "00011111101000000000000000000011";
                        f_reg(361) <= "00100000000111010000000000111100";
                        f_reg(362) <= "00010000000000000000000000000010";
                        f_reg(363) <= "00100000000111010000000000000000";
                        f_reg(364) <= "00010101001101110000000000101110";
                        f_reg(365) <= "10101111101010010000011110110100";
                        f_reg(366) <= "10001100000111010000100000001100";
                        f_reg(367) <= "00011111101000000000000000000011";
                        f_reg(368) <= "00100000000111010000000000111100";
                        f_reg(369) <= "00010000000000000000000000000010";
                        f_reg(370) <= "00100000000111010000000000000000";
                        f_reg(371) <= "00010101010110000000000000100111";
                        f_reg(372) <= "10101111101010100000011110111000";
                        f_reg(373) <= "10001100000111010000100000001100";
                        f_reg(374) <= "00011111101000000000000000000011";
                        f_reg(375) <= "00100000000111010000000000111100";
                        f_reg(376) <= "00010000000000000000000000000010";
                        f_reg(377) <= "00100000000111010000000000000000";
                        f_reg(378) <= "00010101011110010000000000100000";
                        f_reg(379) <= "10101111101010110000011110111100";
                        f_reg(380) <= "10001100000111010000100000001100";
                        f_reg(381) <= "00011111101000000000000000000011";
                        f_reg(382) <= "00100000000111010000000000111100";
                        f_reg(383) <= "00010000000000000000000000000010";
                        f_reg(384) <= "00100000000111010000000000000000";
                        f_reg(385) <= "00010101100110100000000000011001";
                        f_reg(386) <= "10101111101011000000011111000000";
                        f_reg(387) <= "10001100000111010000100000001100";
                        f_reg(388) <= "00011111101000000000000000000011";
                        f_reg(389) <= "00100000000111010000000000111100";
                        f_reg(390) <= "00010000000000000000000000000010";
                        f_reg(391) <= "00100000000111010000000000000000";
                        f_reg(392) <= "00010101101110110000000000010010";
                        f_reg(393) <= "10101111101011010000011111000100";
                        f_reg(394) <= "10001100000111010000100000001100";
                        f_reg(395) <= "00011111101000000000000000000011";
                        f_reg(396) <= "00100000000111010000000000111100";
                        f_reg(397) <= "00010000000000000000000000000010";
                        f_reg(398) <= "00100000000111010000000000000000";
                        f_reg(399) <= "00010101110111000000000000001011";
                        f_reg(400) <= "10101111101011100000011111001000";
                        f_reg(401) <= "10001100000111010000100000001100";
                        f_reg(402) <= "00011111101000000000000000000011";
                        f_reg(403) <= "00100000000111010000000000111100";
                        f_reg(404) <= "00010000000000000000000000000010";
                        f_reg(405) <= "00100000000111010000000000000000";
                        f_reg(406) <= "00010111110111110000000000000100";
                        f_reg(407) <= "10101111101111100000011111001100";
                        f_reg(408) <= "10101100000111010000100000001100";
                        f_reg(409) <= "00010000000000001111111110000100";
                        f_reg(410) <= "10001100000111010000100000001100";
                        f_reg(411) <= "10001111101000010000011110010100";
                        f_reg(412) <= "10001100000111010000100000001100";
                        f_reg(413) <= "10001111101011110000011110010100";
                        f_reg(414) <= "00010100001011111111111111111100";
                        f_reg(415) <= "10001100000111010000100000001100";
                        f_reg(416) <= "10001111101000100000011110011000";
                        f_reg(417) <= "10001100000111010000100000001100";
                        f_reg(418) <= "10001111101100000000011110011000";
                        f_reg(419) <= "00010100010100001111111111111100";
                        f_reg(420) <= "10001100000111010000100000001100";
                        f_reg(421) <= "10001111101000110000011110011100";
                        f_reg(422) <= "10001100000111010000100000001100";
                        f_reg(423) <= "10001111101100010000011110011100";
                        f_reg(424) <= "00010100011100011111111111111100";
                        f_reg(425) <= "10001100000111010000100000001100";
                        f_reg(426) <= "10001111101001000000011110100000";
                        f_reg(427) <= "10001100000111010000100000001100";
                        f_reg(428) <= "10001111101100100000011110100000";
                        f_reg(429) <= "00010100100100101111111111111100";
                        f_reg(430) <= "10001100000111010000100000001100";
                        f_reg(431) <= "10001111101001010000011110100100";
                        f_reg(432) <= "10001100000111010000100000001100";
                        f_reg(433) <= "10001111101100110000011110100100";
                        f_reg(434) <= "00010100101100111111111111111100";
                        f_reg(435) <= "10001100000111010000100000001100";
                        f_reg(436) <= "10001111101001100000011110101000";
                        f_reg(437) <= "10001100000111010000100000001100";
                        f_reg(438) <= "10001111101101000000011110101000";
                        f_reg(439) <= "00010100110101001111111111111100";
                        f_reg(440) <= "10001100000111010000100000001100";
                        f_reg(441) <= "10001111101001110000011110101100";
                        f_reg(442) <= "10001100000111010000100000001100";
                        f_reg(443) <= "10001111101101010000011110101100";
                        f_reg(444) <= "00010100111101011111111111111100";
                        f_reg(445) <= "10001100000111010000100000001100";
                        f_reg(446) <= "10001111101010000000011110110000";
                        f_reg(447) <= "10001100000111010000100000001100";
                        f_reg(448) <= "10001111101101100000011110110000";
                        f_reg(449) <= "00010101000101101111111111111100";
                        f_reg(450) <= "10001100000111010000100000001100";
                        f_reg(451) <= "10001111101010010000011110110100";
                        f_reg(452) <= "10001100000111010000100000001100";
                        f_reg(453) <= "10001111101101110000011110110100";
                        f_reg(454) <= "00010101001101111111111111111100";
                        f_reg(455) <= "10001100000111010000100000001100";
                        f_reg(456) <= "10001111101010100000011110111000";
                        f_reg(457) <= "10001100000111010000100000001100";
                        f_reg(458) <= "10001111101110000000011110111000";
                        f_reg(459) <= "00010101010110001111111111111100";
                        f_reg(460) <= "10001100000111010000100000001100";
                        f_reg(461) <= "10001111101010110000011110111100";
                        f_reg(462) <= "10001100000111010000100000001100";
                        f_reg(463) <= "10001111101110010000011110111100";
                        f_reg(464) <= "00010101011110011111111111111100";
                        f_reg(465) <= "10001100000111010000100000001100";
                        f_reg(466) <= "10001111101011000000011111000000";
                        f_reg(467) <= "10001100000111010000100000001100";
                        f_reg(468) <= "10001111101110100000011111000000";
                        f_reg(469) <= "00010101100110101111111111111100";
                        f_reg(470) <= "10001100000111010000100000001100";
                        f_reg(471) <= "10001111101011010000011111000100";
                        f_reg(472) <= "10001100000111010000100000001100";
                        f_reg(473) <= "10001111101110110000011111000100";
                        f_reg(474) <= "00010101101110111111111111111100";
                        f_reg(475) <= "10001100000111010000100000001100";
                        f_reg(476) <= "10001111101011100000011111001000";
                        f_reg(477) <= "10001100000111010000100000001100";
                        f_reg(478) <= "10001111101111000000011111001000";
                        f_reg(479) <= "00010101110111001111111111111100";
                        f_reg(480) <= "10001100000111010000100000001100";
                        f_reg(481) <= "10001111101111100000011111001100";
                        f_reg(482) <= "10001100000111010000100000001100";
                        f_reg(483) <= "10001111101111110000011111001100";
                        f_reg(484) <= "00010111110111111111111111111100";
                        f_reg(485) <= "00010000000000001111111100111000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000001111100111";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011010100100111011";
                        f_reg(4) <= "00000000000000010001000001000000";
                        f_reg(5) <= "00000000001000000001100000100010";
                        f_reg(6) <= "00000000000000000010010101000010";
                        f_reg(7) <= "00000000011000010010100000000100";
                        f_reg(8) <= "00000000011000110011000000100011";
                        f_reg(9) <= "00000000000000010011100000000110";
                        f_reg(10) <= "00101100101010001111110110000111";
                        f_reg(11) <= "00000000111010000100100000100111";
                        f_reg(12) <= "00100000000010100101111010111001";
                        f_reg(13) <= "00000000000000000000000000000000";
                        f_reg(14) <= "00000001001001100101100000100111";
                        f_reg(15) <= "00000001011000010110000000100110";
                        f_reg(16) <= "00000000000000110110100000100111";
                        f_reg(17) <= "00111001000011101111011001100010";
                        f_reg(18) <= "10101100000011100000010010000100";
                        f_reg(19) <= "00110001100011110110000100110011";
                        f_reg(20) <= "00000000010010101000000000100110";
                        f_reg(21) <= "00000001111100001000100000000110";
                        f_reg(22) <= "00000001111000011001000000100110";
                        f_reg(23) <= "00000000000011001001101111000010";
                        f_reg(24) <= "00000000110100000011000000000110";
                        f_reg(25) <= "00000000101010001010000000100101";
                        f_reg(26) <= "00000010010100111010100000000100";
                        f_reg(27) <= "00000001111001011011000000100001";
                        f_reg(28) <= "00000000000001001011100011000011";
                        f_reg(29) <= "00000010100010011100000000100101";
                        f_reg(30) <= "00000010010100011100100000100010";
                        f_reg(31) <= "00000010111101001101000000100011";
                        f_reg(32) <= "00000001101101101101100000100111";
                        f_reg(33) <= "00000000110110111110000000101010";
                        f_reg(34) <= "00000010000011101110100000100101";
                        f_reg(35) <= "00110100110111101101101111000001";
                        f_reg(36) <= "00000011000110000011100000101010";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00111100000010110110000100010000";
                        f_reg(39) <= "00000000100010110001000000100000";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "00111100000011001110101111111011";
                        f_reg(42) <= "00000000000110000100010010000011";
                        f_reg(43) <= "00000011101101010010100000101010";
                        f_reg(44) <= "00000011100101010100100000100000";
                        f_reg(45) <= "00111001000100011001011011100101";
                        f_reg(46) <= "00000000001011111010000000100001";
                        f_reg(47) <= "00000000000000000000000000000000";
                        f_reg(48) <= "00000000111110100110100000100110";
                        f_reg(49) <= "10101100000001110000010010001000";
                        f_reg(50) <= "00000011001101001011000000100101";
                        f_reg(51) <= "00000011100100011101100000000100";
                        f_reg(52) <= "00000010010010011000000000101011";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00110000101011101011101000001011";
                        f_reg(55) <= "00000000000011000010001000000000";
                        f_reg(56) <= "00000011011011100101100000100000";
                        f_reg(57) <= "00000010110101101100000000100101";
                        f_reg(58) <= "10101100000100110000010010001100";
                        f_reg(59) <= "00000000000000000000000000000000";
                        f_reg(60) <= "10101100000001100000010010010000";
                        f_reg(61) <= "00000000000110001110100000100010";
                        f_reg(62) <= "00000010111010101010100000100001";
                        f_reg(63) <= "00000000100111010100000000000100";
                        f_reg(64) <= "00000001000111100000100000000100";
                        f_reg(65) <= "00101100010011110000110011111111";
                        f_reg(66) <= "00000000000011011101000110000010";
                        f_reg(67) <= "00000000000000010011100111000010";
                        f_reg(68) <= "00000000011101011100100000101010";
                        f_reg(69) <= "00000000111100001010000000101011";
                        f_reg(70) <= "00000000000110011000111110000011";
                        f_reg(71) <= "00000001111100011110000000100010";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "00101101011100101100001010010100";
                        f_reg(74) <= "10101100000111000000010010010100";
                        f_reg(75) <= "10101100000100100000010010011000";
                        f_reg(76) <= "00000000000000000000000000000000";
                        f_reg(77) <= "00110010100010010100000010101111";
                        f_reg(78) <= "00000000000000000000000000000000";
                        f_reg(79) <= "10101100000110100000010010011100";
                        f_reg(80) <= "10101100000010010000010010100000";
                        f_reg(81) <= "00100011111111111111111111111111";
                        f_reg(82) <= "00011111111000001111111110110001";
                        f_reg(83) <= "00010000000000000000000111010100";
                        f_reg(84) <= "00111100000111100000001111100111";
                        f_reg(85) <= "00111100000111110000001111100111";
                        f_reg(86) <= "00000000000111101111010000000010";
                        f_reg(87) <= "00000000000111111111110000000010";
                        f_reg(88) <= "00111100000000011010100100111011";
                        f_reg(89) <= "00111100000011111010100100111011";
                        f_reg(90) <= "00000000000000010001000001000000";
                        f_reg(91) <= "00000000000011111000000001000000";
                        f_reg(92) <= "00000000001000000001100000100010";
                        f_reg(93) <= "00000001111000001000100000100010";
                        f_reg(94) <= "00000000000000000010010101000010";
                        f_reg(95) <= "00000000000000001001010101000010";
                        f_reg(96) <= "00000000011000010010100000000100";
                        f_reg(97) <= "00000010001011111001100000000100";
                        f_reg(98) <= "00000000011000110011000000100011";
                        f_reg(99) <= "00000010001100011010000000100011";
                        f_reg(100) <= "00000000000000010011100000000110";
                        f_reg(101) <= "00000000000011111010100000000110";
                        f_reg(102) <= "00101100101010001111110110000111";
                        f_reg(103) <= "00101110011101101111110110000111";
                        f_reg(104) <= "00000000111010000100100000100111";
                        f_reg(105) <= "00000010101101101011100000100111";
                        f_reg(106) <= "00100000000010100101111010111001";
                        f_reg(107) <= "00100000000110000101111010111001";
                        f_reg(108) <= "00000000000000000000000000000000";
                        f_reg(109) <= "00000000000000000000000000000000";
                        f_reg(110) <= "00000001001001100101100000100111";
                        f_reg(111) <= "00000010111101001100100000100111";
                        f_reg(112) <= "00000001011000010110000000100110";
                        f_reg(113) <= "00000011001011111101000000100110";
                        f_reg(114) <= "00000000000000110110100000100111";
                        f_reg(115) <= "00000000000100011101100000100111";
                        f_reg(116) <= "00111001000011101111011001100010";
                        f_reg(117) <= "00111010110111001111011001100010";
                        f_reg(118) <= "00010101110111000000000100100100";
                        f_reg(119) <= "10101100000011100000010010000100";
                        f_reg(120) <= "00110001100001110110000100110011";
                        f_reg(121) <= "00110011010101010110000100110011";
                        f_reg(122) <= "00000000010010100101100000100110";
                        f_reg(123) <= "00000010000110001100100000100110";
                        f_reg(124) <= "00000000111010110001000000000110";
                        f_reg(125) <= "00000010101110011000000000000110";
                        f_reg(126) <= "00010100011100010000000100011100";
                        f_reg(127) <= "10101100000000110000010010100100";
                        f_reg(128) <= "00000000111000010001100000100110";
                        f_reg(129) <= "00000010101011111000100000100110";
                        f_reg(130) <= "00010101010110000000000100011000";
                        f_reg(131) <= "10101100000010100000010010101000";
                        f_reg(132) <= "00000000000011000101001111000010";
                        f_reg(133) <= "00000000000110101100001111000010";
                        f_reg(134) <= "00000000110010110011000000000110";
                        f_reg(135) <= "00000010100110011010000000000110";
                        f_reg(136) <= "00000000101010000110000000100101";
                        f_reg(137) <= "00000010011101101101000000100101";
                        f_reg(138) <= "00000000011010100100000000000100";
                        f_reg(139) <= "00000010001110001011000000000100";
                        f_reg(140) <= "00010100110101000000000100001110";
                        f_reg(141) <= "10101100000001100000010010101100";
                        f_reg(142) <= "00000000111001010011000000100001";
                        f_reg(143) <= "00000010101100111010000000100001";
                        f_reg(144) <= "00000000000001000010100011000011";
                        f_reg(145) <= "00000000000100101001100011000011";
                        f_reg(146) <= "00010100101100110000000100001000";
                        f_reg(147) <= "10101100000001010000010010110000";
                        f_reg(148) <= "00000001100010010010100000100101";
                        f_reg(149) <= "00000011010101111001100000100101";
                        f_reg(150) <= "00000000011000100100100000100010";
                        f_reg(151) <= "00000010001100001011100000100010";
                        f_reg(152) <= "10001100000000100000010010110000";
                        f_reg(153) <= "10001100000100000000010010110000";
                        f_reg(154) <= "00010100010100001111111111111110";
                        f_reg(155) <= "00010101010110000000000011111111";
                        f_reg(156) <= "10101100000010100000010010110000";
                        f_reg(157) <= "00000000010011000101000000100011";
                        f_reg(158) <= "00000010000110101100000000100011";
                        f_reg(159) <= "00000001101001100110000000100111";
                        f_reg(160) <= "00000011011101001101000000100111";
                        f_reg(161) <= "10001100000011010000010010101100";
                        f_reg(162) <= "10001100000110110000010010101100";
                        f_reg(163) <= "00010101101110111111111111111110";
                        f_reg(164) <= "00000001101011000011000000101010";
                        f_reg(165) <= "00000011011110101010000000101010";
                        f_reg(166) <= "00000001011011100110000000100101";
                        f_reg(167) <= "00000011001111001101000000100101";
                        f_reg(168) <= "00110101101010111101101111000001";
                        f_reg(169) <= "00110111011110011101101111000001";
                        f_reg(170) <= "00000000101001010111000000101010";
                        f_reg(171) <= "00000010011100111110000000101010";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00000000000000000000000000000000";
                        f_reg(174) <= "00010101011110010000000011101100";
                        f_reg(175) <= "10101100000010110000010010101100";
                        f_reg(176) <= "00111100000010110110000100010000";
                        f_reg(177) <= "00111100000110010110000100010000";
                        f_reg(178) <= "00010100010100000000000011101000";
                        f_reg(179) <= "10101100000000100000010010110100";
                        f_reg(180) <= "00000000100010110001000000100000";
                        f_reg(181) <= "00000010010110011000000000100000";
                        f_reg(182) <= "00000000000000000000000000000000";
                        f_reg(183) <= "00000000000000000000000000000000";
                        f_reg(184) <= "00111100000001001110101111111011";
                        f_reg(185) <= "00111100000100101110101111111011";
                        f_reg(186) <= "00000000000001010101110010000011";
                        f_reg(187) <= "00000000000100111100110010000011";
                        f_reg(188) <= "00000001100010000010100000101010";
                        f_reg(189) <= "00000011010101101001100000101010";
                        f_reg(190) <= "00000000110010000110000000100000";
                        f_reg(191) <= "00000010100101101101000000100000";
                        f_reg(192) <= "00111001011010001001011011100101";
                        f_reg(193) <= "00111011001101101001011011100101";
                        f_reg(194) <= "00000000001001110101100000100001";
                        f_reg(195) <= "00000001111101011100100000100001";
                        f_reg(196) <= "00000000000000000000000000000000";
                        f_reg(197) <= "00000000000000000000000000000000";
                        f_reg(198) <= "00000001110010100000100000100110";
                        f_reg(199) <= "00000011100110000111100000100110";
                        f_reg(200) <= "00010101110111000000000011010010";
                        f_reg(201) <= "10101100000011100000010010001000";
                        f_reg(202) <= "00000001001010110011100000100101";
                        f_reg(203) <= "00000010111110011010100000100101";
                        f_reg(204) <= "00000000110010000101000000000100";
                        f_reg(205) <= "00000010100101101100000000000100";
                        f_reg(206) <= "00000000011011000111000000101011";
                        f_reg(207) <= "00000010001110101110000000101011";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00110000101010011011101000001011";
                        f_reg(211) <= "00110010011101111011101000001011";
                        f_reg(212) <= "00000000000001000101101000000000";
                        f_reg(213) <= "00000000000100101100101000000000";
                        f_reg(214) <= "00000001010010010100000000100000";
                        f_reg(215) <= "00000011000101111011000000100000";
                        f_reg(216) <= "00000000111001110011000000100101";
                        f_reg(217) <= "00000010101101011010000000100101";
                        f_reg(218) <= "10001100000000110000010010110000";
                        f_reg(219) <= "10001100000100010000010010110000";
                        f_reg(220) <= "00010100011100011111111111111110";
                        f_reg(221) <= "00010100011100010000000010111101";
                        f_reg(222) <= "10101100000000110000010010001100";
                        f_reg(223) <= "00000000000000000000000000000000";
                        f_reg(224) <= "00000000000000000000000000000000";
                        f_reg(225) <= "00010101101110110000000010111001";
                        f_reg(226) <= "10101100000011010000010010010000";
                        f_reg(227) <= "00000000000001100110000000100010";
                        f_reg(228) <= "00000000000101001101000000100010";
                        f_reg(229) <= "10001100000001010000010010110100";
                        f_reg(230) <= "10001100000100110000010010110100";
                        f_reg(231) <= "00010100101100111111111111111110";
                        f_reg(232) <= "10001100000001000000010010101000";
                        f_reg(233) <= "10001100000100100000010010101000";
                        f_reg(234) <= "00010100100100101111111111111110";
                        f_reg(235) <= "00000000101001000101000000100001";
                        f_reg(236) <= "00000010011100101100000000100001";
                        f_reg(237) <= "00000001011011000100100000000100";
                        f_reg(238) <= "00000011001110101011100000000100";
                        f_reg(239) <= "10001100000001110000010010101100";
                        f_reg(240) <= "10001100000101010000010010101100";
                        f_reg(241) <= "00010100111101011111111111111110";
                        f_reg(242) <= "00000001001001110001100000000100";
                        f_reg(243) <= "00000010111101011000100000000100";
                        f_reg(244) <= "00101100010011010000110011111111";
                        f_reg(245) <= "00101110000110110000110011111111";
                        f_reg(246) <= "00000000000000010011000110000010";
                        f_reg(247) <= "00000000000011111010000110000010";
                        f_reg(248) <= "00000000000000110010100111000010";
                        f_reg(249) <= "00000000000100011001100111000010";
                        f_reg(250) <= "10001100000001000000010010100100";
                        f_reg(251) <= "10001100000100100000010010100100";
                        f_reg(252) <= "00010100100100101111111111111110";
                        f_reg(253) <= "00000000100010100110000000101010";
                        f_reg(254) <= "00000010010110001101000000101010";
                        f_reg(255) <= "00000000101011100101100000101011";
                        f_reg(256) <= "00000010011111001100100000101011";
                        f_reg(257) <= "00000000000011000011111110000011";
                        f_reg(258) <= "00000000000110101010111110000011";
                        f_reg(259) <= "00000001101001110100100000100010";
                        f_reg(260) <= "00000011011101011011100000100010";
                        f_reg(261) <= "00000000000000000000000000000000";
                        f_reg(262) <= "00000000000000000000000000000000";
                        f_reg(263) <= "00101101000000101100001010010100";
                        f_reg(264) <= "00101110110100001100001010010100";
                        f_reg(265) <= "00010101001101110000000010010001";
                        f_reg(266) <= "10101100000010010000010010010100";
                        f_reg(267) <= "00010100010100000000000010001111";
                        f_reg(268) <= "10101100000000100000010010011000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00110001011000010100000010101111";
                        f_reg(272) <= "00110011001011110100000010101111";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00010100110101000000000010000111";
                        f_reg(276) <= "10101100000001100000010010011100";
                        f_reg(277) <= "00010100001011110000000010000101";
                        f_reg(278) <= "10101100000000010000010010100000";
                        f_reg(279) <= "00100011110111011111111100000110";
                        f_reg(280) <= "00010011101000000000000000010111";
                        f_reg(281) <= "00100011110111011111111000001100";
                        f_reg(282) <= "00010011101000000000000000010101";
                        f_reg(283) <= "00100011110111011111110100010010";
                        f_reg(284) <= "00010011101000000000000000010011";
                        f_reg(285) <= "00100011110111101111111111111111";
                        f_reg(286) <= "00100011111111111111111111111111";
                        f_reg(287) <= "00010111110111110000000001111011";
                        f_reg(288) <= "00011111111000001111111100111000";
                        f_reg(289) <= "00010000000000000000000100000110";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "00000000000000000000000000000000";
                        f_reg(293) <= "00000000000000000000000000000000";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "10001100000111010000100000001100";
                        f_reg(304) <= "00011111101000000000000000000011";
                        f_reg(305) <= "00100000000111010000000000111100";
                        f_reg(306) <= "00010000000000000000000000000010";
                        f_reg(307) <= "00100000000111010000000000000000";
                        f_reg(308) <= "00010100001011110000000001100110";
                        f_reg(309) <= "10101111101000010000011110010100";
                        f_reg(310) <= "10001100000111010000100000001100";
                        f_reg(311) <= "00011111101000000000000000000011";
                        f_reg(312) <= "00100000000111010000000000111100";
                        f_reg(313) <= "00010000000000000000000000000010";
                        f_reg(314) <= "00100000000111010000000000000000";
                        f_reg(315) <= "00010100010100000000000001011111";
                        f_reg(316) <= "10101111101000100000011110011000";
                        f_reg(317) <= "10001100000111010000100000001100";
                        f_reg(318) <= "00011111101000000000000000000011";
                        f_reg(319) <= "00100000000111010000000000111100";
                        f_reg(320) <= "00010000000000000000000000000010";
                        f_reg(321) <= "00100000000111010000000000000000";
                        f_reg(322) <= "00010100011100010000000001011000";
                        f_reg(323) <= "10101111101000110000011110011100";
                        f_reg(324) <= "10001100000111010000100000001100";
                        f_reg(325) <= "00011111101000000000000000000011";
                        f_reg(326) <= "00100000000111010000000000111100";
                        f_reg(327) <= "00010000000000000000000000000010";
                        f_reg(328) <= "00100000000111010000000000000000";
                        f_reg(329) <= "00010100100100100000000001010001";
                        f_reg(330) <= "10101111101001000000011110100000";
                        f_reg(331) <= "10001100000111010000100000001100";
                        f_reg(332) <= "00011111101000000000000000000011";
                        f_reg(333) <= "00100000000111010000000000111100";
                        f_reg(334) <= "00010000000000000000000000000010";
                        f_reg(335) <= "00100000000111010000000000000000";
                        f_reg(336) <= "00010100101100110000000001001010";
                        f_reg(337) <= "10101111101001010000011110100100";
                        f_reg(338) <= "10001100000111010000100000001100";
                        f_reg(339) <= "00011111101000000000000000000011";
                        f_reg(340) <= "00100000000111010000000000111100";
                        f_reg(341) <= "00010000000000000000000000000010";
                        f_reg(342) <= "00100000000111010000000000000000";
                        f_reg(343) <= "00010100110101000000000001000011";
                        f_reg(344) <= "10101111101001100000011110101000";
                        f_reg(345) <= "10001100000111010000100000001100";
                        f_reg(346) <= "00011111101000000000000000000011";
                        f_reg(347) <= "00100000000111010000000000111100";
                        f_reg(348) <= "00010000000000000000000000000010";
                        f_reg(349) <= "00100000000111010000000000000000";
                        f_reg(350) <= "00010100111101010000000000111100";
                        f_reg(351) <= "10101111101001110000011110101100";
                        f_reg(352) <= "10001100000111010000100000001100";
                        f_reg(353) <= "00011111101000000000000000000011";
                        f_reg(354) <= "00100000000111010000000000111100";
                        f_reg(355) <= "00010000000000000000000000000010";
                        f_reg(356) <= "00100000000111010000000000000000";
                        f_reg(357) <= "00010101000101100000000000110101";
                        f_reg(358) <= "10101111101010000000011110110000";
                        f_reg(359) <= "10001100000111010000100000001100";
                        f_reg(360) <= "00011111101000000000000000000011";
                        f_reg(361) <= "00100000000111010000000000111100";
                        f_reg(362) <= "00010000000000000000000000000010";
                        f_reg(363) <= "00100000000111010000000000000000";
                        f_reg(364) <= "00010101001101110000000000101110";
                        f_reg(365) <= "10101111101010010000011110110100";
                        f_reg(366) <= "10001100000111010000100000001100";
                        f_reg(367) <= "00011111101000000000000000000011";
                        f_reg(368) <= "00100000000111010000000000111100";
                        f_reg(369) <= "00010000000000000000000000000010";
                        f_reg(370) <= "00100000000111010000000000000000";
                        f_reg(371) <= "00010101010110000000000000100111";
                        f_reg(372) <= "10101111101010100000011110111000";
                        f_reg(373) <= "10001100000111010000100000001100";
                        f_reg(374) <= "00011111101000000000000000000011";
                        f_reg(375) <= "00100000000111010000000000111100";
                        f_reg(376) <= "00010000000000000000000000000010";
                        f_reg(377) <= "00100000000111010000000000000000";
                        f_reg(378) <= "00010101011110010000000000100000";
                        f_reg(379) <= "10101111101010110000011110111100";
                        f_reg(380) <= "10001100000111010000100000001100";
                        f_reg(381) <= "00011111101000000000000000000011";
                        f_reg(382) <= "00100000000111010000000000111100";
                        f_reg(383) <= "00010000000000000000000000000010";
                        f_reg(384) <= "00100000000111010000000000000000";
                        f_reg(385) <= "00010101100110100000000000011001";
                        f_reg(386) <= "10101111101011000000011111000000";
                        f_reg(387) <= "10001100000111010000100000001100";
                        f_reg(388) <= "00011111101000000000000000000011";
                        f_reg(389) <= "00100000000111010000000000111100";
                        f_reg(390) <= "00010000000000000000000000000010";
                        f_reg(391) <= "00100000000111010000000000000000";
                        f_reg(392) <= "00010101101110110000000000010010";
                        f_reg(393) <= "10101111101011010000011111000100";
                        f_reg(394) <= "10001100000111010000100000001100";
                        f_reg(395) <= "00011111101000000000000000000011";
                        f_reg(396) <= "00100000000111010000000000111100";
                        f_reg(397) <= "00010000000000000000000000000010";
                        f_reg(398) <= "00100000000111010000000000000000";
                        f_reg(399) <= "00010101110111000000000000001011";
                        f_reg(400) <= "10101111101011100000011111001000";
                        f_reg(401) <= "10001100000111010000100000001100";
                        f_reg(402) <= "00011111101000000000000000000011";
                        f_reg(403) <= "00100000000111010000000000111100";
                        f_reg(404) <= "00010000000000000000000000000010";
                        f_reg(405) <= "00100000000111010000000000000000";
                        f_reg(406) <= "00010111110111110000000000000100";
                        f_reg(407) <= "10101111101111100000011111001100";
                        f_reg(408) <= "10101100000111010000100000001100";
                        f_reg(409) <= "00010000000000001111111110000100";
                        f_reg(410) <= "10001100000111010000100000001100";
                        f_reg(411) <= "10001111101000010000011110010100";
                        f_reg(412) <= "10001100000111010000100000001100";
                        f_reg(413) <= "10001111101011110000011110010100";
                        f_reg(414) <= "00010100001011111111111111111100";
                        f_reg(415) <= "10001100000111010000100000001100";
                        f_reg(416) <= "10001111101000100000011110011000";
                        f_reg(417) <= "10001100000111010000100000001100";
                        f_reg(418) <= "10001111101100000000011110011000";
                        f_reg(419) <= "00010100010100001111111111111100";
                        f_reg(420) <= "10001100000111010000100000001100";
                        f_reg(421) <= "10001111101000110000011110011100";
                        f_reg(422) <= "10001100000111010000100000001100";
                        f_reg(423) <= "10001111101100010000011110011100";
                        f_reg(424) <= "00010100011100011111111111111100";
                        f_reg(425) <= "10001100000111010000100000001100";
                        f_reg(426) <= "10001111101001000000011110100000";
                        f_reg(427) <= "10001100000111010000100000001100";
                        f_reg(428) <= "10001111101100100000011110100000";
                        f_reg(429) <= "00010100100100101111111111111100";
                        f_reg(430) <= "10001100000111010000100000001100";
                        f_reg(431) <= "10001111101001010000011110100100";
                        f_reg(432) <= "10001100000111010000100000001100";
                        f_reg(433) <= "10001111101100110000011110100100";
                        f_reg(434) <= "00010100101100111111111111111100";
                        f_reg(435) <= "10001100000111010000100000001100";
                        f_reg(436) <= "10001111101001100000011110101000";
                        f_reg(437) <= "10001100000111010000100000001100";
                        f_reg(438) <= "10001111101101000000011110101000";
                        f_reg(439) <= "00010100110101001111111111111100";
                        f_reg(440) <= "10001100000111010000100000001100";
                        f_reg(441) <= "10001111101001110000011110101100";
                        f_reg(442) <= "10001100000111010000100000001100";
                        f_reg(443) <= "10001111101101010000011110101100";
                        f_reg(444) <= "00010100111101011111111111111100";
                        f_reg(445) <= "10001100000111010000100000001100";
                        f_reg(446) <= "10001111101010000000011110110000";
                        f_reg(447) <= "10001100000111010000100000001100";
                        f_reg(448) <= "10001111101101100000011110110000";
                        f_reg(449) <= "00010101000101101111111111111100";
                        f_reg(450) <= "10001100000111010000100000001100";
                        f_reg(451) <= "10001111101010010000011110110100";
                        f_reg(452) <= "10001100000111010000100000001100";
                        f_reg(453) <= "10001111101101110000011110110100";
                        f_reg(454) <= "00010101001101111111111111111100";
                        f_reg(455) <= "10001100000111010000100000001100";
                        f_reg(456) <= "10001111101010100000011110111000";
                        f_reg(457) <= "10001100000111010000100000001100";
                        f_reg(458) <= "10001111101110000000011110111000";
                        f_reg(459) <= "00010101010110001111111111111100";
                        f_reg(460) <= "10001100000111010000100000001100";
                        f_reg(461) <= "10001111101010110000011110111100";
                        f_reg(462) <= "10001100000111010000100000001100";
                        f_reg(463) <= "10001111101110010000011110111100";
                        f_reg(464) <= "00010101011110011111111111111100";
                        f_reg(465) <= "10001100000111010000100000001100";
                        f_reg(466) <= "10001111101011000000011111000000";
                        f_reg(467) <= "10001100000111010000100000001100";
                        f_reg(468) <= "10001111101110100000011111000000";
                        f_reg(469) <= "00010101100110101111111111111100";
                        f_reg(470) <= "10001100000111010000100000001100";
                        f_reg(471) <= "10001111101011010000011111000100";
                        f_reg(472) <= "10001100000111010000100000001100";
                        f_reg(473) <= "10001111101110110000011111000100";
                        f_reg(474) <= "00010101101110111111111111111100";
                        f_reg(475) <= "10001100000111010000100000001100";
                        f_reg(476) <= "10001111101011100000011111001000";
                        f_reg(477) <= "10001100000111010000100000001100";
                        f_reg(478) <= "10001111101111000000011111001000";
                        f_reg(479) <= "00010101110111001111111111111100";
                        f_reg(480) <= "10001100000111010000100000001100";
                        f_reg(481) <= "10001111101111100000011111001100";
                        f_reg(482) <= "10001100000111010000100000001100";
                        f_reg(483) <= "10001111101111110000011111001100";
                        f_reg(484) <= "00010111110111111111111111111100";
                        f_reg(485) <= "00010000000000001111111100111000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000001111100111";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 -22213
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SLL R2 R1 1
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SUB R3 R1 R0
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SRL R4 R0 21
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SLLV R5 R1 R3
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- SUBU R6 R3 R3
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- SRLV R7 R1 R0
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- SLTIU R8 R5 -633
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- NOR R9 R7 R8
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- ADDI R10 R0 24249
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- NOP
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- NOR R11 R9 R6
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- XOR R12 R11 R1
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- NOR R13 R0 R3
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- XORI R14 R8 -2462
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- SW R14 R0 1156
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- ANDI R15 R12 24883
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- XOR R16 R2 R10
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SRLV R17 R16 R15
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- XOR R18 R15 R1
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- SRL R19 R12 15
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- SRLV R6 R16 R6
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- OR R20 R5 R8
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- SLLV R21 R19 R18
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- ADDU R22 R15 R5
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- SRA R23 R4 3
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- OR R24 R20 R9
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- SUB R25 R18 R17
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- SUBU R26 R23 R20
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- NOR R27 R13 R22
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- SLT R28 R6 R27
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- OR R29 R16 R14
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- ORI R30 R6 -9279
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- SLT R7 R24 R24
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- NOP
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- LUI R11 24848
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- ADD R2 R4 R11
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- NOP
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- LUI R12 -5125
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- SRA R8 R24 18
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SLT R5 R29 R21
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- ADD R9 R28 R21
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- XORI R17 R8 -26907
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- ADDU R20 R1 R15
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- NOP
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- XOR R13 R7 R26
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- SW R7 R0 1160
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- OR R22 R25 R20
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SLLV R27 R17 R28
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- SLTU R16 R18 R9
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- NOP
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- ANDI R14 R5 -17909
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SLL R4 R12 8
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- ADD R11 R27 R14
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- OR R24 R22 R22
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- SW R19 R0 1164
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- NOP
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SW R6 R0 1168
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- SUB R29 R0 R24
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- ADDU R21 R23 R10
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- SLLV R8 R29 R4
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- SLLV R1 R30 R8
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- SLTIU R15 R2 3327
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- SRL R26 R13 6
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- SRL R7 R1 7
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- SLT R25 R3 R21
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- SLTU R20 R7 R16
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SRA R17 R25 30
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- SUB R28 R15 R17
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- NOP
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SLTIU R18 R11 -15724
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- SW R28 R0 1172
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- SW R18 R0 1176
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- NOP
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- ANDI R9 R20 16559
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- NOP
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- SW R26 R0 1180
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- SW R9 R0 1184
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- ADDI R31 R31 -1
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- BGTZ R31 -79
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- BEQ R0 R0 468
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- LUI R30 999
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- LUI R31 999
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- SRL R30 R30 16
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SRL R31 R31 16
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- LUI R1 -22213
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- LUI R15 -22213
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- SLL R2 R1 1
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- SLL R16 R15 1
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- SUB R3 R1 R0
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- SUB R17 R15 R0
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- SRL R4 R0 21
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- SRL R18 R0 21
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- SLLV R5 R1 R3
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SLLV R19 R15 R17
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SUBU R6 R3 R3
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- SUBU R20 R17 R17
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- SRLV R7 R1 R0
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- SRLV R21 R15 R0
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- SLTIU R8 R5 -633
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SLTIU R22 R19 -633
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- NOR R9 R7 R8
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- NOR R23 R21 R22
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- ADDI R10 R0 24249
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- ADDI R24 R0 24249
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- NOP
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- NOP
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- NOR R11 R9 R6
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- NOR R25 R23 R20
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- XOR R12 R11 R1
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- XOR R26 R25 R15
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- NOR R13 R0 R3
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- NOR R27 R0 R17
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- XORI R14 R8 -2462
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- XORI R28 R22 -2462
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- BNE R14 R28 292
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- SW R14 R0 1156
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- ANDI R7 R12 24883
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- ANDI R21 R26 24883
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- XOR R11 R2 R10
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- XOR R25 R16 R24
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SRLV R2 R11 R7
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- SRLV R16 R25 R21
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- BNE R3 R17 284
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- SW R3 R0 1188
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- XOR R3 R7 R1
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- XOR R17 R21 R15
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- BNE R10 R24 280
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- SW R10 R0 1192
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- SRL R10 R12 15
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- SRL R24 R26 15
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- SRLV R6 R11 R6
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- SRLV R20 R25 R20
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- OR R12 R5 R8
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- OR R26 R19 R22
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SLLV R8 R10 R3
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- SLLV R22 R24 R17
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- BNE R6 R20 270
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- SW R6 R0 1196
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- ADDU R6 R7 R5
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- ADDU R20 R21 R19
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- SRA R5 R4 3
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- SRA R19 R18 3
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- BNE R5 R19 264
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- SW R5 R0 1200
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- OR R5 R12 R9
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- OR R19 R26 R23
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- SUB R9 R3 R2
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- SUB R23 R17 R16
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- LW R2 R0 1200
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- LW R16 R0 1200
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- BNE R2 R16 -2
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- BNE R10 R24 255
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- SW R10 R0 1200
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- SUBU R10 R2 R12
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- SUBU R24 R16 R26
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- NOR R12 R13 R6
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- NOR R26 R27 R20
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- LW R13 R0 1196
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- LW R27 R0 1196
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- BNE R13 R27 -2
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- SLT R6 R13 R12
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- SLT R20 R27 R26
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- OR R12 R11 R14
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- OR R26 R25 R28
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- ORI R11 R13 -9279
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- ORI R25 R27 -9279
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- SLT R14 R5 R5
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- SLT R28 R19 R19
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- NOP
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- NOP
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- BNE R11 R25 236
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- SW R11 R0 1196
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- LUI R11 24848
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- LUI R25 24848
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- BNE R2 R16 232
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- SW R2 R0 1204
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- ADD R2 R4 R11
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- ADD R16 R18 R25
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- NOP
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- NOP
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- LUI R4 -5125
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- LUI R18 -5125
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- SRA R11 R5 18
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- SRA R25 R19 18
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- SLT R5 R12 R8
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- SLT R19 R26 R22
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- ADD R12 R6 R8
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- ADD R26 R20 R22
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- XORI R8 R11 -26907
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- XORI R22 R25 -26907
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- ADDU R11 R1 R7
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- ADDU R25 R15 R21
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- NOP
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- NOP
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- XOR R1 R14 R10
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- XOR R15 R28 R24
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- BNE R14 R28 210
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- SW R14 R0 1160
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- OR R7 R9 R11
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- OR R21 R23 R25
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- SLLV R10 R8 R6
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- SLLV R24 R22 R20
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- SLTU R14 R3 R12
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- SLTU R28 R17 R26
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- NOP
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- NOP
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- ANDI R9 R5 -17909
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- ANDI R23 R19 -17909
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- SLL R11 R4 8
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- SLL R25 R18 8
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- ADD R8 R10 R9
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- ADD R22 R24 R23
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- OR R6 R7 R7
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- OR R20 R21 R21
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- LW R3 R0 1200
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- LW R17 R0 1200
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- BNE R3 R17 -2
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- BNE R3 R17 189
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- SW R3 R0 1164
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- NOP
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- NOP
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- BNE R13 R27 185
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- SW R13 R0 1168
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- SUB R12 R0 R6
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- SUB R26 R0 R20
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- LW R5 R0 1204
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- LW R19 R0 1204
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- BNE R5 R19 -2
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- LW R4 R0 1192
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- LW R18 R0 1192
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- BNE R4 R18 -2
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- ADDU R10 R5 R4
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- ADDU R24 R19 R18
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- SLLV R9 R12 R11
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- SLLV R23 R26 R25
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- LW R7 R0 1196
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- LW R21 R0 1196
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- BNE R7 R21 -2
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- SLLV R3 R7 R9
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- SLLV R17 R21 R23
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- SLTIU R13 R2 3327
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- SLTIU R27 R16 3327
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- SRL R6 R1 6
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- SRL R20 R15 6
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- SRL R5 R3 7
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- SRL R19 R17 7
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- LW R4 R0 1188
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- LW R18 R0 1188
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- BNE R4 R18 -2
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- SLT R12 R4 R10
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- SLT R26 R18 R24
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- SLTU R11 R5 R14
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- SLTU R25 R19 R28
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- SRA R7 R12 30
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- SRA R21 R26 30
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- SUB R9 R13 R7
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- SUB R23 R27 R21
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- NOP
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- NOP
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- SLTIU R2 R8 -15724
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- SLTIU R16 R22 -15724
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- BNE R9 R23 145
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- SW R9 R0 1172
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- BNE R2 R16 143
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- SW R2 R0 1176
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- NOP
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- NOP
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- ANDI R1 R11 16559
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- ANDI R15 R25 16559
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- NOP
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- NOP
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- BNE R6 R20 135
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- SW R6 R0 1180
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- BNE R1 R15 133
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- SW R1 R0 1184
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- ADDI R29 R30 -250
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- BEQ R29 R0 23
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- ADDI R29 R30 -500
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- BEQ R29 R0 21
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- ADDI R29 R30 -750
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- BEQ R29 R0 19
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- ADDI R30 R30 -1
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- ADDI R31 R31 -1
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- BNE R30 R31 123
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- BGTZ R31 -200
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- BEQ R0 R0 262
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- NOP
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- NOP
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- NOP
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- NOP
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- NOP
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- NOP
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- NOP
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- NOP
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- NOP
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- NOP
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- NOP
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- NOP
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- NOP
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- LW R29 R0 2060
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- BGTZ R29 3
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- ADDI R29 R0 60
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- BEQ R0 R0 2
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- ADDI R29 R0 0
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- BNE R1 R15 102
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- SW R1 R29 1940
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- LW R29 R0 2060
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- BGTZ R29 3
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- ADDI R29 R0 60
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- BEQ R0 R0 2
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- ADDI R29 R0 0
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- BNE R2 R16 95
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- SW R2 R29 1944
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- LW R29 R0 2060
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- BGTZ R29 3
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- ADDI R29 R0 60
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- BEQ R0 R0 2
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- ADDI R29 R0 0
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- BNE R3 R17 88
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- SW R3 R29 1948
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- LW R29 R0 2060
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- BGTZ R29 3
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- ADDI R29 R0 60
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- BEQ R0 R0 2
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- ADDI R29 R0 0
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- BNE R4 R18 81
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- SW R4 R29 1952
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- LW R29 R0 2060
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- BGTZ R29 3
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- ADDI R29 R0 60
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- BEQ R0 R0 2
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- ADDI R29 R0 0
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- BNE R5 R19 74
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- SW R5 R29 1956
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- LW R29 R0 2060
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- BGTZ R29 3
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- ADDI R29 R0 60
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- BEQ R0 R0 2
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- ADDI R29 R0 0
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- BNE R6 R20 67
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- SW R6 R29 1960
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- LW R29 R0 2060
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- BGTZ R29 3
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- ADDI R29 R0 60
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- BEQ R0 R0 2
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- ADDI R29 R0 0
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- BNE R7 R21 60
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- SW R7 R29 1964
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- LW R29 R0 2060
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- BGTZ R29 3
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- ADDI R29 R0 60
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- BEQ R0 R0 2
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- ADDI R29 R0 0
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- BNE R8 R22 53
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- SW R8 R29 1968
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- LW R29 R0 2060
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- BGTZ R29 3
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- ADDI R29 R0 60
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- BEQ R0 R0 2
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- ADDI R29 R0 0
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- BNE R9 R23 46
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- SW R9 R29 1972
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- LW R29 R0 2060
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- BGTZ R29 3
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- ADDI R29 R0 60
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- BEQ R0 R0 2
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- ADDI R29 R0 0
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- BNE R10 R24 39
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- SW R10 R29 1976
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- LW R29 R0 2060
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- BGTZ R29 3
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- ADDI R29 R0 60
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- BEQ R0 R0 2
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- ADDI R29 R0 0
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- BNE R11 R25 32
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- SW R11 R29 1980
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- LW R29 R0 2060
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- BGTZ R29 3
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- ADDI R29 R0 60
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- BEQ R0 R0 2
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- ADDI R29 R0 0
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- BNE R12 R26 25
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- SW R12 R29 1984
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- LW R29 R0 2060
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- BGTZ R29 3
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- ADDI R29 R0 60
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- BEQ R0 R0 2
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- ADDI R29 R0 0
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- BNE R13 R27 18
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- SW R13 R29 1988
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- LW R29 R0 2060
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- BGTZ R29 3
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- ADDI R29 R0 60
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- BEQ R0 R0 2
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- ADDI R29 R0 0
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- BNE R14 R28 11
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- SW R14 R29 1992
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- LW R29 R0 2060
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- BGTZ R29 3
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- ADDI R29 R0 60
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- BEQ R0 R0 2
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- ADDI R29 R0 0
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- BNE R30 R31 4
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- SW R30 R29 1996
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- SW R29 R0 2060
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- BEQ R0 R0 -124
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- LW R29 R0 2060
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- LW R1 R29 1940
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- LW R29 R0 2060
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- LW R15 R29 1940
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- BNE R1 R15 -4
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- LW R29 R0 2060
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- LW R2 R29 1944
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- LW R29 R0 2060
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- LW R16 R29 1944
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- BNE R2 R16 -4
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- LW R29 R0 2060
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- LW R3 R29 1948
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- LW R29 R0 2060
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- LW R17 R29 1948
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- BNE R3 R17 -4
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R29 R0 2060
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R4 R29 1952
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- LW R29 R0 2060
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- LW R18 R29 1952
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- BNE R4 R18 -4
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- LW R29 R0 2060
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- LW R5 R29 1956
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- LW R29 R0 2060
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- LW R19 R29 1956
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- BNE R5 R19 -4
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- LW R29 R0 2060
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- LW R6 R29 1960
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- LW R29 R0 2060
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- LW R20 R29 1960
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- BNE R6 R20 -4
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- LW R29 R0 2060
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- LW R7 R29 1964
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- LW R29 R0 2060
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- LW R21 R29 1964
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- BNE R7 R21 -4
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- LW R29 R0 2060
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- LW R8 R29 1968
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- LW R29 R0 2060
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- LW R22 R29 1968
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- BNE R8 R22 -4
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- LW R29 R0 2060
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- LW R9 R29 1972
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- LW R29 R0 2060
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- LW R23 R29 1972
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- BNE R9 R23 -4
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- LW R29 R0 2060
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- LW R10 R29 1976
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- LW R29 R0 2060
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- LW R24 R29 1976
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- BNE R10 R24 -4
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- LW R29 R0 2060
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- LW R11 R29 1980
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- LW R29 R0 2060
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- LW R25 R29 1980
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- BNE R11 R25 -4
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- LW R29 R0 2060
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- LW R12 R29 1984
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- LW R29 R0 2060
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- LW R26 R29 1984
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- BNE R12 R26 -4
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- LW R29 R0 2060
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- LW R13 R29 1988
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- LW R29 R0 2060
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- LW R27 R29 1988
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- BNE R13 R27 -4
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- LW R29 R0 2060
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- LW R14 R29 1992
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- LW R29 R0 2060
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- LW R28 R29 1992
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- BNE R14 R28 -4
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- LW R29 R0 2060
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- LW R30 R29 1996
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- LW R29 R0 2060
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- LW R31 R29 1996
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- BNE R30 R31 -4
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- BEQ R0 R0 -200
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- NOP
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- NOP
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- NOP
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- NOP
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- NOP
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- NOP
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- NOP
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- NOP
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- NOP
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- NOP
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- NOP
                        f_reg(496) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(497) =>
                        -- NOP
                        f_reg(497) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(498) =>
                        -- NOP
                        f_reg(498) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(499) =>
                        -- NOP
                        f_reg(499) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(500) =>
                        -- NOP
                        f_reg(500) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(501) =>
                        -- NOP
                        f_reg(501) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(502) =>
                        -- NOP
                        f_reg(502) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(503) =>
                        -- NOP
                        f_reg(503) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(504) =>
                        -- NOP
                        f_reg(504) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(505) =>
                        -- NOP
                        f_reg(505) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(506) =>
                        -- NOP
                        f_reg(506) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(507) =>
                        -- NOP
                        f_reg(507) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(508) =>
                        -- NOP
                        f_reg(508) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(509) =>
                        -- NOP
                        f_reg(509) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(510) =>
                        -- NOP
                        f_reg(510) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(511) =>
                        -- NOP
                        f_reg(511) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(512) =>
                        -- NOP
                        f_reg(512) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(513) =>
                        -- NOP
                        f_reg(513) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(514) =>
                        -- NOP
                        f_reg(514) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(515) =>
                        -- NOP
                        f_reg(515) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(516) =>
                        -- NOP
                        f_reg(516) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(517) =>
                        -- NOP
                        f_reg(517) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(518) =>
                        -- NOP
                        f_reg(518) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(519) =>
                        -- NOP
                        f_reg(519) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(520) =>
                        -- NOP
                        f_reg(520) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(521) =>
                        -- NOP
                        f_reg(521) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(522) =>
                        -- NOP
                        f_reg(522) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(523) =>
                        -- NOP
                        f_reg(523) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(524) =>
                        -- NOP
                        f_reg(524) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(525) =>
                        -- NOP
                        f_reg(525) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(526) =>
                        -- NOP
                        f_reg(526) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(527) =>
                        -- NOP
                        f_reg(527) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(528) =>
                        -- NOP
                        f_reg(528) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(529) =>
                        -- NOP
                        f_reg(529) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(530) =>
                        -- NOP
                        f_reg(530) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(531) =>
                        -- NOP
                        f_reg(531) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(532) =>
                        -- NOP
                        f_reg(532) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(533) =>
                        -- NOP
                        f_reg(533) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(534) =>
                        -- NOP
                        f_reg(534) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(535) =>
                        -- NOP
                        f_reg(535) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(536) =>
                        -- NOP
                        f_reg(536) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(537) =>
                        -- NOP
                        f_reg(537) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(538) =>
                        -- NOP
                        f_reg(538) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(539) =>
                        -- NOP
                        f_reg(539) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(540) =>
                        -- NOP
                        f_reg(540) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(541) =>
                        -- NOP
                        f_reg(541) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(542) =>
                        -- NOP
                        f_reg(542) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(543) =>
                        -- NOP
                        f_reg(543) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(544) =>
                        -- NOP
                        f_reg(544) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(545) =>
                        -- NOP
                        f_reg(545) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(546) =>
                        -- NOP
                        f_reg(546) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(547) =>
                        -- NOP
                        f_reg(547) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(548) =>
                        -- NOP
                        f_reg(548) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(549) =>
                        -- NOP
                        f_reg(549) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(550) =>
                        -- NOP
                        f_reg(550) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(551) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011010100100111011";
                        f_reg(4) <= "00000000000000010001000001000000";
                        f_reg(5) <= "00000000001000000001100000100010";
                        f_reg(6) <= "00000000000000000010010101000010";
                        f_reg(7) <= "00000000011000010010100000000100";
                        f_reg(8) <= "00000000011000110011000000100011";
                        f_reg(9) <= "00000000000000010011100000000110";
                        f_reg(10) <= "00101100101010001111110110000111";
                        f_reg(11) <= "00000000111010000100100000100111";
                        f_reg(12) <= "00100000000010100101111010111001";
                        f_reg(13) <= "00000000000000000000000000000000";
                        f_reg(14) <= "00000001001001100101100000100111";
                        f_reg(15) <= "00000001011000010110000000100110";
                        f_reg(16) <= "00000000000000110110100000100111";
                        f_reg(17) <= "00111001000011101111011001100010";
                        f_reg(18) <= "10101100000011100000010010000100";
                        f_reg(19) <= "00110001100011110110000100110011";
                        f_reg(20) <= "00000000010010101000000000100110";
                        f_reg(21) <= "00000001111100001000100000000110";
                        f_reg(22) <= "00000001111000011001000000100110";
                        f_reg(23) <= "00000000000011001001101111000010";
                        f_reg(24) <= "00000000110100000011000000000110";
                        f_reg(25) <= "00000000101010001010000000100101";
                        f_reg(26) <= "00000010010100111010100000000100";
                        f_reg(27) <= "00000001111001011011000000100001";
                        f_reg(28) <= "00000000000001001011100011000011";
                        f_reg(29) <= "00000010100010011100000000100101";
                        f_reg(30) <= "00000010010100011100100000100010";
                        f_reg(31) <= "00000010111101001101000000100011";
                        f_reg(32) <= "00000001101101101101100000100111";
                        f_reg(33) <= "00000000110110111110000000101010";
                        f_reg(34) <= "00000010000011101110100000100101";
                        f_reg(35) <= "00110100110111101101101111000001";
                        f_reg(36) <= "00000011000110000011100000101010";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00111100000010110110000100010000";
                        f_reg(39) <= "00000000100010110001000000100000";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "00111100000011001110101111111011";
                        f_reg(42) <= "00000000000110000100010010000011";
                        f_reg(43) <= "00000011101101010010100000101010";
                        f_reg(44) <= "00000011100101010100100000100000";
                        f_reg(45) <= "00111001000100011001011011100101";
                        f_reg(46) <= "00000000001011111010000000100001";
                        f_reg(47) <= "00000000000000000000000000000000";
                        f_reg(48) <= "00000000111110100110100000100110";
                        f_reg(49) <= "10101100000001110000010010001000";
                        f_reg(50) <= "00000011001101001011000000100101";
                        f_reg(51) <= "00000011100100011101100000000100";
                        f_reg(52) <= "00000010010010011000000000101011";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00110000101011101011101000001011";
                        f_reg(55) <= "00000000000011000010001000000000";
                        f_reg(56) <= "00000011011011100101100000100000";
                        f_reg(57) <= "00000010110101101100000000100101";
                        f_reg(58) <= "10101100000100110000010010001100";
                        f_reg(59) <= "00000000000000000000000000000000";
                        f_reg(60) <= "10101100000001100000010010010000";
                        f_reg(61) <= "00000000000110001110100000100010";
                        f_reg(62) <= "00000010111010101010100000100001";
                        f_reg(63) <= "00000000100111010100000000000100";
                        f_reg(64) <= "00000001000111100000100000000100";
                        f_reg(65) <= "00101100010011110000110011111111";
                        f_reg(66) <= "00000000000011011101000110000010";
                        f_reg(67) <= "00000000000000010011100111000010";
                        f_reg(68) <= "00000000011101011100100000101010";
                        f_reg(69) <= "00000000111100001010000000101011";
                        f_reg(70) <= "00000000000110011000111110000011";
                        f_reg(71) <= "00000001111100011110000000100010";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "00101101011100101100001010010100";
                        f_reg(74) <= "10101100000111000000010010010100";
                        f_reg(75) <= "10101100000100100000010010011000";
                        f_reg(76) <= "00000000000000000000000000000000";
                        f_reg(77) <= "00110010100010010100000010101111";
                        f_reg(78) <= "00000000000000000000000000000000";
                        f_reg(79) <= "10101100000110100000010010011100";
                        f_reg(80) <= "10101100000010010000010010100000";
                        f_reg(81) <= "00100011111111111111111111111111";
                        f_reg(82) <= "00011111111000001111111110110001";
                        f_reg(83) <= "00010000000000000000000111010100";
                        f_reg(84) <= "00111100000111100000001111100111";
                        f_reg(85) <= "00111100000111110000001111100111";
                        f_reg(86) <= "00000000000111101111010000000010";
                        f_reg(87) <= "00000000000111111111110000000010";
                        f_reg(88) <= "00111100000000011010100100111011";
                        f_reg(89) <= "00111100000011111010100100111011";
                        f_reg(90) <= "00000000000000010001000001000000";
                        f_reg(91) <= "00000000000011111000000001000000";
                        f_reg(92) <= "00000000001000000001100000100010";
                        f_reg(93) <= "00000001111000001000100000100010";
                        f_reg(94) <= "00000000000000000010010101000010";
                        f_reg(95) <= "00000000000000001001010101000010";
                        f_reg(96) <= "00000000011000010010100000000100";
                        f_reg(97) <= "00000010001011111001100000000100";
                        f_reg(98) <= "00000000011000110011000000100011";
                        f_reg(99) <= "00000010001100011010000000100011";
                        f_reg(100) <= "00000000000000010011100000000110";
                        f_reg(101) <= "00000000000011111010100000000110";
                        f_reg(102) <= "00101100101010001111110110000111";
                        f_reg(103) <= "00101110011101101111110110000111";
                        f_reg(104) <= "00000000111010000100100000100111";
                        f_reg(105) <= "00000010101101101011100000100111";
                        f_reg(106) <= "00100000000010100101111010111001";
                        f_reg(107) <= "00100000000110000101111010111001";
                        f_reg(108) <= "00000000000000000000000000000000";
                        f_reg(109) <= "00000000000000000000000000000000";
                        f_reg(110) <= "00000001001001100101100000100111";
                        f_reg(111) <= "00000010111101001100100000100111";
                        f_reg(112) <= "00000001011000010110000000100110";
                        f_reg(113) <= "00000011001011111101000000100110";
                        f_reg(114) <= "00000000000000110110100000100111";
                        f_reg(115) <= "00000000000100011101100000100111";
                        f_reg(116) <= "00111001000011101111011001100010";
                        f_reg(117) <= "00111010110111001111011001100010";
                        f_reg(118) <= "00010101110111000000000100100100";
                        f_reg(119) <= "10101100000011100000010010000100";
                        f_reg(120) <= "00110001100001110110000100110011";
                        f_reg(121) <= "00110011010101010110000100110011";
                        f_reg(122) <= "00000000010010100101100000100110";
                        f_reg(123) <= "00000010000110001100100000100110";
                        f_reg(124) <= "00000000111010110001000000000110";
                        f_reg(125) <= "00000010101110011000000000000110";
                        f_reg(126) <= "00010100011100010000000100011100";
                        f_reg(127) <= "10101100000000110000010010100100";
                        f_reg(128) <= "00000000111000010001100000100110";
                        f_reg(129) <= "00000010101011111000100000100110";
                        f_reg(130) <= "00010101010110000000000100011000";
                        f_reg(131) <= "10101100000010100000010010101000";
                        f_reg(132) <= "00000000000011000101001111000010";
                        f_reg(133) <= "00000000000110101100001111000010";
                        f_reg(134) <= "00000000110010110011000000000110";
                        f_reg(135) <= "00000010100110011010000000000110";
                        f_reg(136) <= "00000000101010000110000000100101";
                        f_reg(137) <= "00000010011101101101000000100101";
                        f_reg(138) <= "00000000011010100100000000000100";
                        f_reg(139) <= "00000010001110001011000000000100";
                        f_reg(140) <= "00010100110101000000000100001110";
                        f_reg(141) <= "10101100000001100000010010101100";
                        f_reg(142) <= "00000000111001010011000000100001";
                        f_reg(143) <= "00000010101100111010000000100001";
                        f_reg(144) <= "00000000000001000010100011000011";
                        f_reg(145) <= "00000000000100101001100011000011";
                        f_reg(146) <= "00010100101100110000000100001000";
                        f_reg(147) <= "10101100000001010000010010110000";
                        f_reg(148) <= "00000001100010010010100000100101";
                        f_reg(149) <= "00000011010101111001100000100101";
                        f_reg(150) <= "00000000011000100100100000100010";
                        f_reg(151) <= "00000010001100001011100000100010";
                        f_reg(152) <= "10001100000000100000010010110000";
                        f_reg(153) <= "10001100000100000000010010110000";
                        f_reg(154) <= "00010100010100001111111111111110";
                        f_reg(155) <= "00010101010110000000000011111111";
                        f_reg(156) <= "10101100000010100000010010110000";
                        f_reg(157) <= "00000000010011000101000000100011";
                        f_reg(158) <= "00000010000110101100000000100011";
                        f_reg(159) <= "00000001101001100110000000100111";
                        f_reg(160) <= "00000011011101001101000000100111";
                        f_reg(161) <= "10001100000011010000010010101100";
                        f_reg(162) <= "10001100000110110000010010101100";
                        f_reg(163) <= "00010101101110111111111111111110";
                        f_reg(164) <= "00000001101011000011000000101010";
                        f_reg(165) <= "00000011011110101010000000101010";
                        f_reg(166) <= "00000001011011100110000000100101";
                        f_reg(167) <= "00000011001111001101000000100101";
                        f_reg(168) <= "00110101101010111101101111000001";
                        f_reg(169) <= "00110111011110011101101111000001";
                        f_reg(170) <= "00000000101001010111000000101010";
                        f_reg(171) <= "00000010011100111110000000101010";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00000000000000000000000000000000";
                        f_reg(174) <= "00010101011110010000000011101100";
                        f_reg(175) <= "10101100000010110000010010101100";
                        f_reg(176) <= "00111100000010110110000100010000";
                        f_reg(177) <= "00111100000110010110000100010000";
                        f_reg(178) <= "00010100010100000000000011101000";
                        f_reg(179) <= "10101100000000100000010010110100";
                        f_reg(180) <= "00000000100010110001000000100000";
                        f_reg(181) <= "00000010010110011000000000100000";
                        f_reg(182) <= "00000000000000000000000000000000";
                        f_reg(183) <= "00000000000000000000000000000000";
                        f_reg(184) <= "00111100000001001110101111111011";
                        f_reg(185) <= "00111100000100101110101111111011";
                        f_reg(186) <= "00000000000001010101110010000011";
                        f_reg(187) <= "00000000000100111100110010000011";
                        f_reg(188) <= "00000001100010000010100000101010";
                        f_reg(189) <= "00000011010101101001100000101010";
                        f_reg(190) <= "00000000110010000110000000100000";
                        f_reg(191) <= "00000010100101101101000000100000";
                        f_reg(192) <= "00111001011010001001011011100101";
                        f_reg(193) <= "00111011001101101001011011100101";
                        f_reg(194) <= "00000000001001110101100000100001";
                        f_reg(195) <= "00000001111101011100100000100001";
                        f_reg(196) <= "00000000000000000000000000000000";
                        f_reg(197) <= "00000000000000000000000000000000";
                        f_reg(198) <= "00000001110010100000100000100110";
                        f_reg(199) <= "00000011100110000111100000100110";
                        f_reg(200) <= "00010101110111000000000011010010";
                        f_reg(201) <= "10101100000011100000010010001000";
                        f_reg(202) <= "00000001001010110011100000100101";
                        f_reg(203) <= "00000010111110011010100000100101";
                        f_reg(204) <= "00000000110010000101000000000100";
                        f_reg(205) <= "00000010100101101100000000000100";
                        f_reg(206) <= "00000000011011000111000000101011";
                        f_reg(207) <= "00000010001110101110000000101011";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00110000101010011011101000001011";
                        f_reg(211) <= "00110010011101111011101000001011";
                        f_reg(212) <= "00000000000001000101101000000000";
                        f_reg(213) <= "00000000000100101100101000000000";
                        f_reg(214) <= "00000001010010010100000000100000";
                        f_reg(215) <= "00000011000101111011000000100000";
                        f_reg(216) <= "00000000111001110011000000100101";
                        f_reg(217) <= "00000010101101011010000000100101";
                        f_reg(218) <= "10001100000000110000010010110000";
                        f_reg(219) <= "10001100000100010000010010110000";
                        f_reg(220) <= "00010100011100011111111111111110";
                        f_reg(221) <= "00010100011100010000000010111101";
                        f_reg(222) <= "10101100000000110000010010001100";
                        f_reg(223) <= "00000000000000000000000000000000";
                        f_reg(224) <= "00000000000000000000000000000000";
                        f_reg(225) <= "00010101101110110000000010111001";
                        f_reg(226) <= "10101100000011010000010010010000";
                        f_reg(227) <= "00000000000001100110000000100010";
                        f_reg(228) <= "00000000000101001101000000100010";
                        f_reg(229) <= "10001100000001010000010010110100";
                        f_reg(230) <= "10001100000100110000010010110100";
                        f_reg(231) <= "00010100101100111111111111111110";
                        f_reg(232) <= "10001100000001000000010010101000";
                        f_reg(233) <= "10001100000100100000010010101000";
                        f_reg(234) <= "00010100100100101111111111111110";
                        f_reg(235) <= "00000000101001000101000000100001";
                        f_reg(236) <= "00000010011100101100000000100001";
                        f_reg(237) <= "00000001011011000100100000000100";
                        f_reg(238) <= "00000011001110101011100000000100";
                        f_reg(239) <= "10001100000001110000010010101100";
                        f_reg(240) <= "10001100000101010000010010101100";
                        f_reg(241) <= "00010100111101011111111111111110";
                        f_reg(242) <= "00000001001001110001100000000100";
                        f_reg(243) <= "00000010111101011000100000000100";
                        f_reg(244) <= "00101100010011010000110011111111";
                        f_reg(245) <= "00101110000110110000110011111111";
                        f_reg(246) <= "00000000000000010011000110000010";
                        f_reg(247) <= "00000000000011111010000110000010";
                        f_reg(248) <= "00000000000000110010100111000010";
                        f_reg(249) <= "00000000000100011001100111000010";
                        f_reg(250) <= "10001100000001000000010010100100";
                        f_reg(251) <= "10001100000100100000010010100100";
                        f_reg(252) <= "00010100100100101111111111111110";
                        f_reg(253) <= "00000000100010100110000000101010";
                        f_reg(254) <= "00000010010110001101000000101010";
                        f_reg(255) <= "00000000101011100101100000101011";
                        f_reg(256) <= "00000010011111001100100000101011";
                        f_reg(257) <= "00000000000011000011111110000011";
                        f_reg(258) <= "00000000000110101010111110000011";
                        f_reg(259) <= "00000001101001110100100000100010";
                        f_reg(260) <= "00000011011101011011100000100010";
                        f_reg(261) <= "00000000000000000000000000000000";
                        f_reg(262) <= "00000000000000000000000000000000";
                        f_reg(263) <= "00101101000000101100001010010100";
                        f_reg(264) <= "00101110110100001100001010010100";
                        f_reg(265) <= "00010101001101110000000010010001";
                        f_reg(266) <= "10101100000010010000010010010100";
                        f_reg(267) <= "00010100010100000000000010001111";
                        f_reg(268) <= "10101100000000100000010010011000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00110001011000010100000010101111";
                        f_reg(272) <= "00110011001011110100000010101111";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00010100110101000000000010000111";
                        f_reg(276) <= "10101100000001100000010010011100";
                        f_reg(277) <= "00010100001011110000000010000101";
                        f_reg(278) <= "10101100000000010000010010100000";
                        f_reg(279) <= "00100011110111011111111100000110";
                        f_reg(280) <= "00010011101000000000000000010111";
                        f_reg(281) <= "00100011110111011111111000001100";
                        f_reg(282) <= "00010011101000000000000000010101";
                        f_reg(283) <= "00100011110111011111110100010010";
                        f_reg(284) <= "00010011101000000000000000010011";
                        f_reg(285) <= "00100011110111101111111111111111";
                        f_reg(286) <= "00100011111111111111111111111111";
                        f_reg(287) <= "00010111110111110000000001111011";
                        f_reg(288) <= "00011111111000001111111100111000";
                        f_reg(289) <= "00010000000000000000000100000110";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "00000000000000000000000000000000";
                        f_reg(293) <= "00000000000000000000000000000000";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "10001100000111010000100000001100";
                        f_reg(304) <= "00011111101000000000000000000011";
                        f_reg(305) <= "00100000000111010000000000111100";
                        f_reg(306) <= "00010000000000000000000000000010";
                        f_reg(307) <= "00100000000111010000000000000000";
                        f_reg(308) <= "00010100001011110000000001100110";
                        f_reg(309) <= "10101111101000010000011110010100";
                        f_reg(310) <= "10001100000111010000100000001100";
                        f_reg(311) <= "00011111101000000000000000000011";
                        f_reg(312) <= "00100000000111010000000000111100";
                        f_reg(313) <= "00010000000000000000000000000010";
                        f_reg(314) <= "00100000000111010000000000000000";
                        f_reg(315) <= "00010100010100000000000001011111";
                        f_reg(316) <= "10101111101000100000011110011000";
                        f_reg(317) <= "10001100000111010000100000001100";
                        f_reg(318) <= "00011111101000000000000000000011";
                        f_reg(319) <= "00100000000111010000000000111100";
                        f_reg(320) <= "00010000000000000000000000000010";
                        f_reg(321) <= "00100000000111010000000000000000";
                        f_reg(322) <= "00010100011100010000000001011000";
                        f_reg(323) <= "10101111101000110000011110011100";
                        f_reg(324) <= "10001100000111010000100000001100";
                        f_reg(325) <= "00011111101000000000000000000011";
                        f_reg(326) <= "00100000000111010000000000111100";
                        f_reg(327) <= "00010000000000000000000000000010";
                        f_reg(328) <= "00100000000111010000000000000000";
                        f_reg(329) <= "00010100100100100000000001010001";
                        f_reg(330) <= "10101111101001000000011110100000";
                        f_reg(331) <= "10001100000111010000100000001100";
                        f_reg(332) <= "00011111101000000000000000000011";
                        f_reg(333) <= "00100000000111010000000000111100";
                        f_reg(334) <= "00010000000000000000000000000010";
                        f_reg(335) <= "00100000000111010000000000000000";
                        f_reg(336) <= "00010100101100110000000001001010";
                        f_reg(337) <= "10101111101001010000011110100100";
                        f_reg(338) <= "10001100000111010000100000001100";
                        f_reg(339) <= "00011111101000000000000000000011";
                        f_reg(340) <= "00100000000111010000000000111100";
                        f_reg(341) <= "00010000000000000000000000000010";
                        f_reg(342) <= "00100000000111010000000000000000";
                        f_reg(343) <= "00010100110101000000000001000011";
                        f_reg(344) <= "10101111101001100000011110101000";
                        f_reg(345) <= "10001100000111010000100000001100";
                        f_reg(346) <= "00011111101000000000000000000011";
                        f_reg(347) <= "00100000000111010000000000111100";
                        f_reg(348) <= "00010000000000000000000000000010";
                        f_reg(349) <= "00100000000111010000000000000000";
                        f_reg(350) <= "00010100111101010000000000111100";
                        f_reg(351) <= "10101111101001110000011110101100";
                        f_reg(352) <= "10001100000111010000100000001100";
                        f_reg(353) <= "00011111101000000000000000000011";
                        f_reg(354) <= "00100000000111010000000000111100";
                        f_reg(355) <= "00010000000000000000000000000010";
                        f_reg(356) <= "00100000000111010000000000000000";
                        f_reg(357) <= "00010101000101100000000000110101";
                        f_reg(358) <= "10101111101010000000011110110000";
                        f_reg(359) <= "10001100000111010000100000001100";
                        f_reg(360) <= "00011111101000000000000000000011";
                        f_reg(361) <= "00100000000111010000000000111100";
                        f_reg(362) <= "00010000000000000000000000000010";
                        f_reg(363) <= "00100000000111010000000000000000";
                        f_reg(364) <= "00010101001101110000000000101110";
                        f_reg(365) <= "10101111101010010000011110110100";
                        f_reg(366) <= "10001100000111010000100000001100";
                        f_reg(367) <= "00011111101000000000000000000011";
                        f_reg(368) <= "00100000000111010000000000111100";
                        f_reg(369) <= "00010000000000000000000000000010";
                        f_reg(370) <= "00100000000111010000000000000000";
                        f_reg(371) <= "00010101010110000000000000100111";
                        f_reg(372) <= "10101111101010100000011110111000";
                        f_reg(373) <= "10001100000111010000100000001100";
                        f_reg(374) <= "00011111101000000000000000000011";
                        f_reg(375) <= "00100000000111010000000000111100";
                        f_reg(376) <= "00010000000000000000000000000010";
                        f_reg(377) <= "00100000000111010000000000000000";
                        f_reg(378) <= "00010101011110010000000000100000";
                        f_reg(379) <= "10101111101010110000011110111100";
                        f_reg(380) <= "10001100000111010000100000001100";
                        f_reg(381) <= "00011111101000000000000000000011";
                        f_reg(382) <= "00100000000111010000000000111100";
                        f_reg(383) <= "00010000000000000000000000000010";
                        f_reg(384) <= "00100000000111010000000000000000";
                        f_reg(385) <= "00010101100110100000000000011001";
                        f_reg(386) <= "10101111101011000000011111000000";
                        f_reg(387) <= "10001100000111010000100000001100";
                        f_reg(388) <= "00011111101000000000000000000011";
                        f_reg(389) <= "00100000000111010000000000111100";
                        f_reg(390) <= "00010000000000000000000000000010";
                        f_reg(391) <= "00100000000111010000000000000000";
                        f_reg(392) <= "00010101101110110000000000010010";
                        f_reg(393) <= "10101111101011010000011111000100";
                        f_reg(394) <= "10001100000111010000100000001100";
                        f_reg(395) <= "00011111101000000000000000000011";
                        f_reg(396) <= "00100000000111010000000000111100";
                        f_reg(397) <= "00010000000000000000000000000010";
                        f_reg(398) <= "00100000000111010000000000000000";
                        f_reg(399) <= "00010101110111000000000000001011";
                        f_reg(400) <= "10101111101011100000011111001000";
                        f_reg(401) <= "10001100000111010000100000001100";
                        f_reg(402) <= "00011111101000000000000000000011";
                        f_reg(403) <= "00100000000111010000000000111100";
                        f_reg(404) <= "00010000000000000000000000000010";
                        f_reg(405) <= "00100000000111010000000000000000";
                        f_reg(406) <= "00010111110111110000000000000100";
                        f_reg(407) <= "10101111101111100000011111001100";
                        f_reg(408) <= "10101100000111010000100000001100";
                        f_reg(409) <= "00010000000000001111111110000100";
                        f_reg(410) <= "10001100000111010000100000001100";
                        f_reg(411) <= "10001111101000010000011110010100";
                        f_reg(412) <= "10001100000111010000100000001100";
                        f_reg(413) <= "10001111101011110000011110010100";
                        f_reg(414) <= "00010100001011111111111111111100";
                        f_reg(415) <= "10001100000111010000100000001100";
                        f_reg(416) <= "10001111101000100000011110011000";
                        f_reg(417) <= "10001100000111010000100000001100";
                        f_reg(418) <= "10001111101100000000011110011000";
                        f_reg(419) <= "00010100010100001111111111111100";
                        f_reg(420) <= "10001100000111010000100000001100";
                        f_reg(421) <= "10001111101000110000011110011100";
                        f_reg(422) <= "10001100000111010000100000001100";
                        f_reg(423) <= "10001111101100010000011110011100";
                        f_reg(424) <= "00010100011100011111111111111100";
                        f_reg(425) <= "10001100000111010000100000001100";
                        f_reg(426) <= "10001111101001000000011110100000";
                        f_reg(427) <= "10001100000111010000100000001100";
                        f_reg(428) <= "10001111101100100000011110100000";
                        f_reg(429) <= "00010100100100101111111111111100";
                        f_reg(430) <= "10001100000111010000100000001100";
                        f_reg(431) <= "10001111101001010000011110100100";
                        f_reg(432) <= "10001100000111010000100000001100";
                        f_reg(433) <= "10001111101100110000011110100100";
                        f_reg(434) <= "00010100101100111111111111111100";
                        f_reg(435) <= "10001100000111010000100000001100";
                        f_reg(436) <= "10001111101001100000011110101000";
                        f_reg(437) <= "10001100000111010000100000001100";
                        f_reg(438) <= "10001111101101000000011110101000";
                        f_reg(439) <= "00010100110101001111111111111100";
                        f_reg(440) <= "10001100000111010000100000001100";
                        f_reg(441) <= "10001111101001110000011110101100";
                        f_reg(442) <= "10001100000111010000100000001100";
                        f_reg(443) <= "10001111101101010000011110101100";
                        f_reg(444) <= "00010100111101011111111111111100";
                        f_reg(445) <= "10001100000111010000100000001100";
                        f_reg(446) <= "10001111101010000000011110110000";
                        f_reg(447) <= "10001100000111010000100000001100";
                        f_reg(448) <= "10001111101101100000011110110000";
                        f_reg(449) <= "00010101000101101111111111111100";
                        f_reg(450) <= "10001100000111010000100000001100";
                        f_reg(451) <= "10001111101010010000011110110100";
                        f_reg(452) <= "10001100000111010000100000001100";
                        f_reg(453) <= "10001111101101110000011110110100";
                        f_reg(454) <= "00010101001101111111111111111100";
                        f_reg(455) <= "10001100000111010000100000001100";
                        f_reg(456) <= "10001111101010100000011110111000";
                        f_reg(457) <= "10001100000111010000100000001100";
                        f_reg(458) <= "10001111101110000000011110111000";
                        f_reg(459) <= "00010101010110001111111111111100";
                        f_reg(460) <= "10001100000111010000100000001100";
                        f_reg(461) <= "10001111101010110000011110111100";
                        f_reg(462) <= "10001100000111010000100000001100";
                        f_reg(463) <= "10001111101110010000011110111100";
                        f_reg(464) <= "00010101011110011111111111111100";
                        f_reg(465) <= "10001100000111010000100000001100";
                        f_reg(466) <= "10001111101011000000011111000000";
                        f_reg(467) <= "10001100000111010000100000001100";
                        f_reg(468) <= "10001111101110100000011111000000";
                        f_reg(469) <= "00010101100110101111111111111100";
                        f_reg(470) <= "10001100000111010000100000001100";
                        f_reg(471) <= "10001111101011010000011111000100";
                        f_reg(472) <= "10001100000111010000100000001100";
                        f_reg(473) <= "10001111101110110000011111000100";
                        f_reg(474) <= "00010101101110111111111111111100";
                        f_reg(475) <= "10001100000111010000100000001100";
                        f_reg(476) <= "10001111101011100000011111001000";
                        f_reg(477) <= "10001100000111010000100000001100";
                        f_reg(478) <= "10001111101111000000011111001000";
                        f_reg(479) <= "00010101110111001111111111111100";
                        f_reg(480) <= "10001100000111010000100000001100";
                        f_reg(481) <= "10001111101111100000011111001100";
                        f_reg(482) <= "10001100000111010000100000001100";
                        f_reg(483) <= "10001111101111110000011111001100";
                        f_reg(484) <= "00010111110111111111111111111100";
                        f_reg(485) <= "00010000000000001111111100111000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000001111100111";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011010100100111011";
                        f_reg(4) <= "00000000000000010001000001000000";
                        f_reg(5) <= "00000000001000000001100000100010";
                        f_reg(6) <= "00000000000000000010010101000010";
                        f_reg(7) <= "00000000011000010010100000000100";
                        f_reg(8) <= "00000000011000110011000000100011";
                        f_reg(9) <= "00000000000000010011100000000110";
                        f_reg(10) <= "00101100101010001111110110000111";
                        f_reg(11) <= "00000000111010000100100000100111";
                        f_reg(12) <= "00100000000010100101111010111001";
                        f_reg(13) <= "00000000000000000000000000000000";
                        f_reg(14) <= "00000001001001100101100000100111";
                        f_reg(15) <= "00000001011000010110000000100110";
                        f_reg(16) <= "00000000000000110110100000100111";
                        f_reg(17) <= "00111001000011101111011001100010";
                        f_reg(18) <= "10101100000011100000010010000100";
                        f_reg(19) <= "00110001100011110110000100110011";
                        f_reg(20) <= "00000000010010101000000000100110";
                        f_reg(21) <= "00000001111100001000100000000110";
                        f_reg(22) <= "00000001111000011001000000100110";
                        f_reg(23) <= "00000000000011001001101111000010";
                        f_reg(24) <= "00000000110100000011000000000110";
                        f_reg(25) <= "00000000101010001010000000100101";
                        f_reg(26) <= "00000010010100111010100000000100";
                        f_reg(27) <= "00000001111001011011000000100001";
                        f_reg(28) <= "00000000000001001011100011000011";
                        f_reg(29) <= "00000010100010011100000000100101";
                        f_reg(30) <= "00000010010100011100100000100010";
                        f_reg(31) <= "00000010111101001101000000100011";
                        f_reg(32) <= "00000001101101101101100000100111";
                        f_reg(33) <= "00000000110110111110000000101010";
                        f_reg(34) <= "00000010000011101110100000100101";
                        f_reg(35) <= "00110100110111101101101111000001";
                        f_reg(36) <= "00000011000110000011100000101010";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00111100000010110110000100010000";
                        f_reg(39) <= "00000000100010110001000000100000";
                        f_reg(40) <= "00000000000000000000000000000000";
                        f_reg(41) <= "00111100000011001110101111111011";
                        f_reg(42) <= "00000000000110000100010010000011";
                        f_reg(43) <= "00000011101101010010100000101010";
                        f_reg(44) <= "00000011100101010100100000100000";
                        f_reg(45) <= "00111001000100011001011011100101";
                        f_reg(46) <= "00000000001011111010000000100001";
                        f_reg(47) <= "00000000000000000000000000000000";
                        f_reg(48) <= "00000000111110100110100000100110";
                        f_reg(49) <= "10101100000001110000010010001000";
                        f_reg(50) <= "00000011001101001011000000100101";
                        f_reg(51) <= "00000011100100011101100000000100";
                        f_reg(52) <= "00000010010010011000000000101011";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00110000101011101011101000001011";
                        f_reg(55) <= "00000000000011000010001000000000";
                        f_reg(56) <= "00000011011011100101100000100000";
                        f_reg(57) <= "00000010110101101100000000100101";
                        f_reg(58) <= "10101100000100110000010010001100";
                        f_reg(59) <= "00000000000000000000000000000000";
                        f_reg(60) <= "10101100000001100000010010010000";
                        f_reg(61) <= "00000000000110001110100000100010";
                        f_reg(62) <= "00000010111010101010100000100001";
                        f_reg(63) <= "00000000100111010100000000000100";
                        f_reg(64) <= "00000001000111100000100000000100";
                        f_reg(65) <= "00101100010011110000110011111111";
                        f_reg(66) <= "00000000000011011101000110000010";
                        f_reg(67) <= "00000000000000010011100111000010";
                        f_reg(68) <= "00000000011101011100100000101010";
                        f_reg(69) <= "00000000111100001010000000101011";
                        f_reg(70) <= "00000000000110011000111110000011";
                        f_reg(71) <= "00000001111100011110000000100010";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "00101101011100101100001010010100";
                        f_reg(74) <= "10101100000111000000010010010100";
                        f_reg(75) <= "10101100000100100000010010011000";
                        f_reg(76) <= "00000000000000000000000000000000";
                        f_reg(77) <= "00110010100010010100000010101111";
                        f_reg(78) <= "00000000000000000000000000000000";
                        f_reg(79) <= "10101100000110100000010010011100";
                        f_reg(80) <= "10101100000010010000010010100000";
                        f_reg(81) <= "00100011111111111111111111111111";
                        f_reg(82) <= "00011111111000001111111110110001";
                        f_reg(83) <= "00010000000000000000000111010100";
                        f_reg(84) <= "00111100000111100000001111100111";
                        f_reg(85) <= "00111100000111110000001111100111";
                        f_reg(86) <= "00000000000111101111010000000010";
                        f_reg(87) <= "00000000000111111111110000000010";
                        f_reg(88) <= "00111100000000011010100100111011";
                        f_reg(89) <= "00111100000011111010100100111011";
                        f_reg(90) <= "00000000000000010001000001000000";
                        f_reg(91) <= "00000000000011111000000001000000";
                        f_reg(92) <= "00000000001000000001100000100010";
                        f_reg(93) <= "00000001111000001000100000100010";
                        f_reg(94) <= "00000000000000000010010101000010";
                        f_reg(95) <= "00000000000000001001010101000010";
                        f_reg(96) <= "00000000011000010010100000000100";
                        f_reg(97) <= "00000010001011111001100000000100";
                        f_reg(98) <= "00000000011000110011000000100011";
                        f_reg(99) <= "00000010001100011010000000100011";
                        f_reg(100) <= "00000000000000010011100000000110";
                        f_reg(101) <= "00000000000011111010100000000110";
                        f_reg(102) <= "00101100101010001111110110000111";
                        f_reg(103) <= "00101110011101101111110110000111";
                        f_reg(104) <= "00000000111010000100100000100111";
                        f_reg(105) <= "00000010101101101011100000100111";
                        f_reg(106) <= "00100000000010100101111010111001";
                        f_reg(107) <= "00100000000110000101111010111001";
                        f_reg(108) <= "00000000000000000000000000000000";
                        f_reg(109) <= "00000000000000000000000000000000";
                        f_reg(110) <= "00000001001001100101100000100111";
                        f_reg(111) <= "00000010111101001100100000100111";
                        f_reg(112) <= "00000001011000010110000000100110";
                        f_reg(113) <= "00000011001011111101000000100110";
                        f_reg(114) <= "00000000000000110110100000100111";
                        f_reg(115) <= "00000000000100011101100000100111";
                        f_reg(116) <= "00111001000011101111011001100010";
                        f_reg(117) <= "00111010110111001111011001100010";
                        f_reg(118) <= "00010101110111000000000100100100";
                        f_reg(119) <= "10101100000011100000010010000100";
                        f_reg(120) <= "00110001100001110110000100110011";
                        f_reg(121) <= "00110011010101010110000100110011";
                        f_reg(122) <= "00000000010010100101100000100110";
                        f_reg(123) <= "00000010000110001100100000100110";
                        f_reg(124) <= "00000000111010110001000000000110";
                        f_reg(125) <= "00000010101110011000000000000110";
                        f_reg(126) <= "00010100011100010000000100011100";
                        f_reg(127) <= "10101100000000110000010010100100";
                        f_reg(128) <= "00000000111000010001100000100110";
                        f_reg(129) <= "00000010101011111000100000100110";
                        f_reg(130) <= "00010101010110000000000100011000";
                        f_reg(131) <= "10101100000010100000010010101000";
                        f_reg(132) <= "00000000000011000101001111000010";
                        f_reg(133) <= "00000000000110101100001111000010";
                        f_reg(134) <= "00000000110010110011000000000110";
                        f_reg(135) <= "00000010100110011010000000000110";
                        f_reg(136) <= "00000000101010000110000000100101";
                        f_reg(137) <= "00000010011101101101000000100101";
                        f_reg(138) <= "00000000011010100100000000000100";
                        f_reg(139) <= "00000010001110001011000000000100";
                        f_reg(140) <= "00010100110101000000000100001110";
                        f_reg(141) <= "10101100000001100000010010101100";
                        f_reg(142) <= "00000000111001010011000000100001";
                        f_reg(143) <= "00000010101100111010000000100001";
                        f_reg(144) <= "00000000000001000010100011000011";
                        f_reg(145) <= "00000000000100101001100011000011";
                        f_reg(146) <= "00010100101100110000000100001000";
                        f_reg(147) <= "10101100000001010000010010110000";
                        f_reg(148) <= "00000001100010010010100000100101";
                        f_reg(149) <= "00000011010101111001100000100101";
                        f_reg(150) <= "00000000011000100100100000100010";
                        f_reg(151) <= "00000010001100001011100000100010";
                        f_reg(152) <= "10001100000000100000010010110000";
                        f_reg(153) <= "10001100000100000000010010110000";
                        f_reg(154) <= "00010100010100001111111111111110";
                        f_reg(155) <= "00010101010110000000000011111111";
                        f_reg(156) <= "10101100000010100000010010110000";
                        f_reg(157) <= "00000000010011000101000000100011";
                        f_reg(158) <= "00000010000110101100000000100011";
                        f_reg(159) <= "00000001101001100110000000100111";
                        f_reg(160) <= "00000011011101001101000000100111";
                        f_reg(161) <= "10001100000011010000010010101100";
                        f_reg(162) <= "10001100000110110000010010101100";
                        f_reg(163) <= "00010101101110111111111111111110";
                        f_reg(164) <= "00000001101011000011000000101010";
                        f_reg(165) <= "00000011011110101010000000101010";
                        f_reg(166) <= "00000001011011100110000000100101";
                        f_reg(167) <= "00000011001111001101000000100101";
                        f_reg(168) <= "00110101101010111101101111000001";
                        f_reg(169) <= "00110111011110011101101111000001";
                        f_reg(170) <= "00000000101001010111000000101010";
                        f_reg(171) <= "00000010011100111110000000101010";
                        f_reg(172) <= "00000000000000000000000000000000";
                        f_reg(173) <= "00000000000000000000000000000000";
                        f_reg(174) <= "00010101011110010000000011101100";
                        f_reg(175) <= "10101100000010110000010010101100";
                        f_reg(176) <= "00111100000010110110000100010000";
                        f_reg(177) <= "00111100000110010110000100010000";
                        f_reg(178) <= "00010100010100000000000011101000";
                        f_reg(179) <= "10101100000000100000010010110100";
                        f_reg(180) <= "00000000100010110001000000100000";
                        f_reg(181) <= "00000010010110011000000000100000";
                        f_reg(182) <= "00000000000000000000000000000000";
                        f_reg(183) <= "00000000000000000000000000000000";
                        f_reg(184) <= "00111100000001001110101111111011";
                        f_reg(185) <= "00111100000100101110101111111011";
                        f_reg(186) <= "00000000000001010101110010000011";
                        f_reg(187) <= "00000000000100111100110010000011";
                        f_reg(188) <= "00000001100010000010100000101010";
                        f_reg(189) <= "00000011010101101001100000101010";
                        f_reg(190) <= "00000000110010000110000000100000";
                        f_reg(191) <= "00000010100101101101000000100000";
                        f_reg(192) <= "00111001011010001001011011100101";
                        f_reg(193) <= "00111011001101101001011011100101";
                        f_reg(194) <= "00000000001001110101100000100001";
                        f_reg(195) <= "00000001111101011100100000100001";
                        f_reg(196) <= "00000000000000000000000000000000";
                        f_reg(197) <= "00000000000000000000000000000000";
                        f_reg(198) <= "00000001110010100000100000100110";
                        f_reg(199) <= "00000011100110000111100000100110";
                        f_reg(200) <= "00010101110111000000000011010010";
                        f_reg(201) <= "10101100000011100000010010001000";
                        f_reg(202) <= "00000001001010110011100000100101";
                        f_reg(203) <= "00000010111110011010100000100101";
                        f_reg(204) <= "00000000110010000101000000000100";
                        f_reg(205) <= "00000010100101101100000000000100";
                        f_reg(206) <= "00000000011011000111000000101011";
                        f_reg(207) <= "00000010001110101110000000101011";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00110000101010011011101000001011";
                        f_reg(211) <= "00110010011101111011101000001011";
                        f_reg(212) <= "00000000000001000101101000000000";
                        f_reg(213) <= "00000000000100101100101000000000";
                        f_reg(214) <= "00000001010010010100000000100000";
                        f_reg(215) <= "00000011000101111011000000100000";
                        f_reg(216) <= "00000000111001110011000000100101";
                        f_reg(217) <= "00000010101101011010000000100101";
                        f_reg(218) <= "10001100000000110000010010110000";
                        f_reg(219) <= "10001100000100010000010010110000";
                        f_reg(220) <= "00010100011100011111111111111110";
                        f_reg(221) <= "00010100011100010000000010111101";
                        f_reg(222) <= "10101100000000110000010010001100";
                        f_reg(223) <= "00000000000000000000000000000000";
                        f_reg(224) <= "00000000000000000000000000000000";
                        f_reg(225) <= "00010101101110110000000010111001";
                        f_reg(226) <= "10101100000011010000010010010000";
                        f_reg(227) <= "00000000000001100110000000100010";
                        f_reg(228) <= "00000000000101001101000000100010";
                        f_reg(229) <= "10001100000001010000010010110100";
                        f_reg(230) <= "10001100000100110000010010110100";
                        f_reg(231) <= "00010100101100111111111111111110";
                        f_reg(232) <= "10001100000001000000010010101000";
                        f_reg(233) <= "10001100000100100000010010101000";
                        f_reg(234) <= "00010100100100101111111111111110";
                        f_reg(235) <= "00000000101001000101000000100001";
                        f_reg(236) <= "00000010011100101100000000100001";
                        f_reg(237) <= "00000001011011000100100000000100";
                        f_reg(238) <= "00000011001110101011100000000100";
                        f_reg(239) <= "10001100000001110000010010101100";
                        f_reg(240) <= "10001100000101010000010010101100";
                        f_reg(241) <= "00010100111101011111111111111110";
                        f_reg(242) <= "00000001001001110001100000000100";
                        f_reg(243) <= "00000010111101011000100000000100";
                        f_reg(244) <= "00101100010011010000110011111111";
                        f_reg(245) <= "00101110000110110000110011111111";
                        f_reg(246) <= "00000000000000010011000110000010";
                        f_reg(247) <= "00000000000011111010000110000010";
                        f_reg(248) <= "00000000000000110010100111000010";
                        f_reg(249) <= "00000000000100011001100111000010";
                        f_reg(250) <= "10001100000001000000010010100100";
                        f_reg(251) <= "10001100000100100000010010100100";
                        f_reg(252) <= "00010100100100101111111111111110";
                        f_reg(253) <= "00000000100010100110000000101010";
                        f_reg(254) <= "00000010010110001101000000101010";
                        f_reg(255) <= "00000000101011100101100000101011";
                        f_reg(256) <= "00000010011111001100100000101011";
                        f_reg(257) <= "00000000000011000011111110000011";
                        f_reg(258) <= "00000000000110101010111110000011";
                        f_reg(259) <= "00000001101001110100100000100010";
                        f_reg(260) <= "00000011011101011011100000100010";
                        f_reg(261) <= "00000000000000000000000000000000";
                        f_reg(262) <= "00000000000000000000000000000000";
                        f_reg(263) <= "00101101000000101100001010010100";
                        f_reg(264) <= "00101110110100001100001010010100";
                        f_reg(265) <= "00010101001101110000000010010001";
                        f_reg(266) <= "10101100000010010000010010010100";
                        f_reg(267) <= "00010100010100000000000010001111";
                        f_reg(268) <= "10101100000000100000010010011000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00110001011000010100000010101111";
                        f_reg(272) <= "00110011001011110100000010101111";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00010100110101000000000010000111";
                        f_reg(276) <= "10101100000001100000010010011100";
                        f_reg(277) <= "00010100001011110000000010000101";
                        f_reg(278) <= "10101100000000010000010010100000";
                        f_reg(279) <= "00100011110111011111111100000110";
                        f_reg(280) <= "00010011101000000000000000010111";
                        f_reg(281) <= "00100011110111011111111000001100";
                        f_reg(282) <= "00010011101000000000000000010101";
                        f_reg(283) <= "00100011110111011111110100010010";
                        f_reg(284) <= "00010011101000000000000000010011";
                        f_reg(285) <= "00100011110111101111111111111111";
                        f_reg(286) <= "00100011111111111111111111111111";
                        f_reg(287) <= "00010111110111110000000001111011";
                        f_reg(288) <= "00011111111000001111111100111000";
                        f_reg(289) <= "00010000000000000000000100000110";
                        f_reg(290) <= "00000000000000000000000000000000";
                        f_reg(291) <= "00000000000000000000000000000000";
                        f_reg(292) <= "00000000000000000000000000000000";
                        f_reg(293) <= "00000000000000000000000000000000";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "10001100000111010000100000001100";
                        f_reg(304) <= "00011111101000000000000000000011";
                        f_reg(305) <= "00100000000111010000000000111100";
                        f_reg(306) <= "00010000000000000000000000000010";
                        f_reg(307) <= "00100000000111010000000000000000";
                        f_reg(308) <= "00010100001011110000000001100110";
                        f_reg(309) <= "10101111101000010000011110010100";
                        f_reg(310) <= "10001100000111010000100000001100";
                        f_reg(311) <= "00011111101000000000000000000011";
                        f_reg(312) <= "00100000000111010000000000111100";
                        f_reg(313) <= "00010000000000000000000000000010";
                        f_reg(314) <= "00100000000111010000000000000000";
                        f_reg(315) <= "00010100010100000000000001011111";
                        f_reg(316) <= "10101111101000100000011110011000";
                        f_reg(317) <= "10001100000111010000100000001100";
                        f_reg(318) <= "00011111101000000000000000000011";
                        f_reg(319) <= "00100000000111010000000000111100";
                        f_reg(320) <= "00010000000000000000000000000010";
                        f_reg(321) <= "00100000000111010000000000000000";
                        f_reg(322) <= "00010100011100010000000001011000";
                        f_reg(323) <= "10101111101000110000011110011100";
                        f_reg(324) <= "10001100000111010000100000001100";
                        f_reg(325) <= "00011111101000000000000000000011";
                        f_reg(326) <= "00100000000111010000000000111100";
                        f_reg(327) <= "00010000000000000000000000000010";
                        f_reg(328) <= "00100000000111010000000000000000";
                        f_reg(329) <= "00010100100100100000000001010001";
                        f_reg(330) <= "10101111101001000000011110100000";
                        f_reg(331) <= "10001100000111010000100000001100";
                        f_reg(332) <= "00011111101000000000000000000011";
                        f_reg(333) <= "00100000000111010000000000111100";
                        f_reg(334) <= "00010000000000000000000000000010";
                        f_reg(335) <= "00100000000111010000000000000000";
                        f_reg(336) <= "00010100101100110000000001001010";
                        f_reg(337) <= "10101111101001010000011110100100";
                        f_reg(338) <= "10001100000111010000100000001100";
                        f_reg(339) <= "00011111101000000000000000000011";
                        f_reg(340) <= "00100000000111010000000000111100";
                        f_reg(341) <= "00010000000000000000000000000010";
                        f_reg(342) <= "00100000000111010000000000000000";
                        f_reg(343) <= "00010100110101000000000001000011";
                        f_reg(344) <= "10101111101001100000011110101000";
                        f_reg(345) <= "10001100000111010000100000001100";
                        f_reg(346) <= "00011111101000000000000000000011";
                        f_reg(347) <= "00100000000111010000000000111100";
                        f_reg(348) <= "00010000000000000000000000000010";
                        f_reg(349) <= "00100000000111010000000000000000";
                        f_reg(350) <= "00010100111101010000000000111100";
                        f_reg(351) <= "10101111101001110000011110101100";
                        f_reg(352) <= "10001100000111010000100000001100";
                        f_reg(353) <= "00011111101000000000000000000011";
                        f_reg(354) <= "00100000000111010000000000111100";
                        f_reg(355) <= "00010000000000000000000000000010";
                        f_reg(356) <= "00100000000111010000000000000000";
                        f_reg(357) <= "00010101000101100000000000110101";
                        f_reg(358) <= "10101111101010000000011110110000";
                        f_reg(359) <= "10001100000111010000100000001100";
                        f_reg(360) <= "00011111101000000000000000000011";
                        f_reg(361) <= "00100000000111010000000000111100";
                        f_reg(362) <= "00010000000000000000000000000010";
                        f_reg(363) <= "00100000000111010000000000000000";
                        f_reg(364) <= "00010101001101110000000000101110";
                        f_reg(365) <= "10101111101010010000011110110100";
                        f_reg(366) <= "10001100000111010000100000001100";
                        f_reg(367) <= "00011111101000000000000000000011";
                        f_reg(368) <= "00100000000111010000000000111100";
                        f_reg(369) <= "00010000000000000000000000000010";
                        f_reg(370) <= "00100000000111010000000000000000";
                        f_reg(371) <= "00010101010110000000000000100111";
                        f_reg(372) <= "10101111101010100000011110111000";
                        f_reg(373) <= "10001100000111010000100000001100";
                        f_reg(374) <= "00011111101000000000000000000011";
                        f_reg(375) <= "00100000000111010000000000111100";
                        f_reg(376) <= "00010000000000000000000000000010";
                        f_reg(377) <= "00100000000111010000000000000000";
                        f_reg(378) <= "00010101011110010000000000100000";
                        f_reg(379) <= "10101111101010110000011110111100";
                        f_reg(380) <= "10001100000111010000100000001100";
                        f_reg(381) <= "00011111101000000000000000000011";
                        f_reg(382) <= "00100000000111010000000000111100";
                        f_reg(383) <= "00010000000000000000000000000010";
                        f_reg(384) <= "00100000000111010000000000000000";
                        f_reg(385) <= "00010101100110100000000000011001";
                        f_reg(386) <= "10101111101011000000011111000000";
                        f_reg(387) <= "10001100000111010000100000001100";
                        f_reg(388) <= "00011111101000000000000000000011";
                        f_reg(389) <= "00100000000111010000000000111100";
                        f_reg(390) <= "00010000000000000000000000000010";
                        f_reg(391) <= "00100000000111010000000000000000";
                        f_reg(392) <= "00010101101110110000000000010010";
                        f_reg(393) <= "10101111101011010000011111000100";
                        f_reg(394) <= "10001100000111010000100000001100";
                        f_reg(395) <= "00011111101000000000000000000011";
                        f_reg(396) <= "00100000000111010000000000111100";
                        f_reg(397) <= "00010000000000000000000000000010";
                        f_reg(398) <= "00100000000111010000000000000000";
                        f_reg(399) <= "00010101110111000000000000001011";
                        f_reg(400) <= "10101111101011100000011111001000";
                        f_reg(401) <= "10001100000111010000100000001100";
                        f_reg(402) <= "00011111101000000000000000000011";
                        f_reg(403) <= "00100000000111010000000000111100";
                        f_reg(404) <= "00010000000000000000000000000010";
                        f_reg(405) <= "00100000000111010000000000000000";
                        f_reg(406) <= "00010111110111110000000000000100";
                        f_reg(407) <= "10101111101111100000011111001100";
                        f_reg(408) <= "10101100000111010000100000001100";
                        f_reg(409) <= "00010000000000001111111110000100";
                        f_reg(410) <= "10001100000111010000100000001100";
                        f_reg(411) <= "10001111101000010000011110010100";
                        f_reg(412) <= "10001100000111010000100000001100";
                        f_reg(413) <= "10001111101011110000011110010100";
                        f_reg(414) <= "00010100001011111111111111111100";
                        f_reg(415) <= "10001100000111010000100000001100";
                        f_reg(416) <= "10001111101000100000011110011000";
                        f_reg(417) <= "10001100000111010000100000001100";
                        f_reg(418) <= "10001111101100000000011110011000";
                        f_reg(419) <= "00010100010100001111111111111100";
                        f_reg(420) <= "10001100000111010000100000001100";
                        f_reg(421) <= "10001111101000110000011110011100";
                        f_reg(422) <= "10001100000111010000100000001100";
                        f_reg(423) <= "10001111101100010000011110011100";
                        f_reg(424) <= "00010100011100011111111111111100";
                        f_reg(425) <= "10001100000111010000100000001100";
                        f_reg(426) <= "10001111101001000000011110100000";
                        f_reg(427) <= "10001100000111010000100000001100";
                        f_reg(428) <= "10001111101100100000011110100000";
                        f_reg(429) <= "00010100100100101111111111111100";
                        f_reg(430) <= "10001100000111010000100000001100";
                        f_reg(431) <= "10001111101001010000011110100100";
                        f_reg(432) <= "10001100000111010000100000001100";
                        f_reg(433) <= "10001111101100110000011110100100";
                        f_reg(434) <= "00010100101100111111111111111100";
                        f_reg(435) <= "10001100000111010000100000001100";
                        f_reg(436) <= "10001111101001100000011110101000";
                        f_reg(437) <= "10001100000111010000100000001100";
                        f_reg(438) <= "10001111101101000000011110101000";
                        f_reg(439) <= "00010100110101001111111111111100";
                        f_reg(440) <= "10001100000111010000100000001100";
                        f_reg(441) <= "10001111101001110000011110101100";
                        f_reg(442) <= "10001100000111010000100000001100";
                        f_reg(443) <= "10001111101101010000011110101100";
                        f_reg(444) <= "00010100111101011111111111111100";
                        f_reg(445) <= "10001100000111010000100000001100";
                        f_reg(446) <= "10001111101010000000011110110000";
                        f_reg(447) <= "10001100000111010000100000001100";
                        f_reg(448) <= "10001111101101100000011110110000";
                        f_reg(449) <= "00010101000101101111111111111100";
                        f_reg(450) <= "10001100000111010000100000001100";
                        f_reg(451) <= "10001111101010010000011110110100";
                        f_reg(452) <= "10001100000111010000100000001100";
                        f_reg(453) <= "10001111101101110000011110110100";
                        f_reg(454) <= "00010101001101111111111111111100";
                        f_reg(455) <= "10001100000111010000100000001100";
                        f_reg(456) <= "10001111101010100000011110111000";
                        f_reg(457) <= "10001100000111010000100000001100";
                        f_reg(458) <= "10001111101110000000011110111000";
                        f_reg(459) <= "00010101010110001111111111111100";
                        f_reg(460) <= "10001100000111010000100000001100";
                        f_reg(461) <= "10001111101010110000011110111100";
                        f_reg(462) <= "10001100000111010000100000001100";
                        f_reg(463) <= "10001111101110010000011110111100";
                        f_reg(464) <= "00010101011110011111111111111100";
                        f_reg(465) <= "10001100000111010000100000001100";
                        f_reg(466) <= "10001111101011000000011111000000";
                        f_reg(467) <= "10001100000111010000100000001100";
                        f_reg(468) <= "10001111101110100000011111000000";
                        f_reg(469) <= "00010101100110101111111111111100";
                        f_reg(470) <= "10001100000111010000100000001100";
                        f_reg(471) <= "10001111101011010000011111000100";
                        f_reg(472) <= "10001100000111010000100000001100";
                        f_reg(473) <= "10001111101110110000011111000100";
                        f_reg(474) <= "00010101101110111111111111111100";
                        f_reg(475) <= "10001100000111010000100000001100";
                        f_reg(476) <= "10001111101011100000011111001000";
                        f_reg(477) <= "10001100000111010000100000001100";
                        f_reg(478) <= "10001111101111000000011111001000";
                        f_reg(479) <= "00010101110111001111111111111100";
                        f_reg(480) <= "10001100000111010000100000001100";
                        f_reg(481) <= "10001111101111100000011111001100";
                        f_reg(482) <= "10001100000111010000100000001100";
                        f_reg(483) <= "10001111101111110000011111001100";
                        f_reg(484) <= "00010111110111111111111111111100";
                        f_reg(485) <= "00010000000000001111111100111000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000001111100111";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test77_Reg_COMBINED;
