--| Test59_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:12:04
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test59_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test59_Reg_COMBINED;

architecture a_Test59_Reg_COMBINED of Test59_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 521) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 521) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100", --  495 - 1980
      "00000000000000000000011111000000", --  496 - 1984
      "00000000000000000000011111000100", --  497 - 1988
      "00000000000000000000011111001000", --  498 - 1992
      "00000000000000000000011111001100", --  499 - 1996
      "00000000000000000000011111010000", --  500 - 2000
      "00000000000000000000011111010100", --  501 - 2004
      "00000000000000000000011111011000", --  502 - 2008
      "00000000000000000000011111011100", --  503 - 2012
      "00000000000000000000011111100000", --  504 - 2016
      "00000000000000000000011111100100", --  505 - 2020
      "00000000000000000000011111101000", --  506 - 2024
      "00000000000000000000011111101100", --  507 - 2028
      "00000000000000000000011111110000", --  508 - 2032
      "00000000000000000000011111110100", --  509 - 2036
      "00000000000000000000011111111000", --  510 - 2040
      "00000000000000000000011111111100", --  511 - 2044
      "00000000000000000000100000000000", --  512 - 2048
      "00000000000000000000100000000100", --  513 - 2052
      "00000000000000000000100000001000", --  514 - 2056
      "00000000000000000000100000001100", --  515 - 2060
      "00000000000000000000100000010000", --  516 - 2064
      "00000000000000000000100000010100", --  517 - 2068
      "00000000000000000000100000011000", --  518 - 2072
      "00000000000000000000100000011100", --  519 - 2076
      "00000000000000000000100000100000");--  520 - 2080

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000011110001011000110", --    2 -    8
      "00000000000000010001000000100011", --    3 -   12
      "00110000010000110010110010110100", --    4 -   16
      "00000000000000100010010111000011", --    5 -   20
      "00000000100000110010100000100101", --    6 -   24
      "00000000101001000011000000100111", --    7 -   28
      "00000000000001000011100000100000", --    8 -   32
      "00000000110001100100000000100110", --    9 -   36
      "00000000011001110100100000000110", --   10 -   40
      "00000000100001010101000000101011", --   11 -   44
      "00111100000010111011000100000110", --   12 -   48
      "00000000001000000110000000100111", --   13 -   52
      "00000000000000000000000000000000", --   14 -   56
      "00000000100010110110100000100001", --   15 -   60
      "00000000100000100111000000100100", --   16 -   64
      "00000001110010010111100000000111", --   17 -   68
      "00000000000010101000010101000011", --   18 -   72
      "00000001110010011000100000100110", --   19 -   76
      "00000001010011011001000000100001", --   20 -   80
      "00111100000100111111100001001000", --   21 -   84
      "00110000100101000010101000100001", --   22 -   88
      "00110010001101011110100101000110", --   23 -   92
      "00000000000001000010010101000011", --   24 -   96
      "00110001011101100000001011101110", --   25 -  100
      "00000001111001111011100000100011", --   26 -  104
      "00000000000000000000000000000000", --   27 -  108
      "00000010000000111100000000100010", --   28 -  112
      "00000010101101111100100000100101", --   29 -  116
      "00000001110100101101000000100111", --   30 -  120
      "00000000101011101101100000100101", --   31 -  124
      "00000011001000111110000000000110", --   32 -  128
      "00110011100111010110101000011011", --   33 -  132
      "00000010101101111111000000100101", --   34 -  136
      "00100011000001101011100111011001", --   35 -  140
      "00000000000100110000110101000011", --   36 -  144
      "00111100000000101011111011010101", --   37 -  148
      "00000001011110110100100000100101", --   38 -  152
      "00000011010000010101000000100000", --   39 -  156
      "00000001010101000110100000100001", --   40 -  160
      "00101101101100010110111101000101", --   41 -  164
      "00000000110111010111100000000111", --   42 -  168
      "00000010010011110011100000100100", --   43 -  172
      "00000000010100011000000000100101", --   44 -  176
      "00000010110100000010100000100110", --   45 -  180
      "00101110110011100011000111001011", --   46 -  184
      "00101001000000111100000010111011", --   47 -  188
      "00000000101001101110000000100001", --   48 -  192
      "00000011011011001010100000100110", --   49 -  196
      "00000010101111101011100000101011", --   50 -  200
      "00000000000000000000000000000000", --   51 -  204
      "00000000111001001100000000000111", --   52 -  208
      "10101100000010000000010000011100", --   53 -  212
      "00000001011011101001100000100110", --   54 -  216
      "00000000000000000000000000000000", --   55 -  220
      "00000000000000111101000111000010", --   56 -  224
      "00000000000111000000111001000011", --   57 -  228
      "00100110111010101001000110111000", --   58 -  232
      "10101100000110010000010000100000", --   59 -  236
      "00110100101101001111111000101001", --   60 -  240
      "00100011010011010010111110011100", --   61 -  244
      "00000001001101001110100000100001", --   62 -  248
      "00000000000000000000000000000000", --   63 -  252
      "00000011000000001001000000101011", --   64 -  256
      "00000011101000010111100000100101", --   65 -  260
      "00000000000000000000000000000000", --   66 -  264
      "00000001010011110001000000100111", --   67 -  268
      "10101100000011010000010000100100", --   68 -  272
      "10101100000100100000010000101000", --   69 -  276
      "10101100000100110000010000101100", --   70 -  280
      "00000000000000000000000000000000", --   71 -  284
      "10101100000000100000010000110000", --   72 -  288
      "00100011111111111111111111111111", --   73 -  292
      "00011111111000001111111110111000", --   74 -  296
      "00010000000000000000000110111101", --   75 -  300
      "00111100000111100000001111100111", --   76 -  304
      "00111100000111110000001111100111", --   77 -  308
      "00000000000111101111010000000010", --   78 -  312
      "00000000000111111111110000000010", --   79 -  316
      "00111100000000011110001011000110", --   80 -  320
      "00111100000011111110001011000110", --   81 -  324
      "00000000000000010001000000100011", --   82 -  328
      "00000000000011111000000000100011", --   83 -  332
      "00110000010000110010110010110100", --   84 -  336
      "00110010000100010010110010110100", --   85 -  340
      "00000000000000100010010111000011", --   86 -  344
      "00000000000100001001010111000011", --   87 -  348
      "00000000100000110010100000100101", --   88 -  352
      "00000010010100011001100000100101", --   89 -  356
      "00000000101001000011000000100111", --   90 -  360
      "00000010011100101010000000100111", --   91 -  364
      "00000000000001000011100000100000", --   92 -  368
      "00000000000100101010100000100000", --   93 -  372
      "00000000110001100100000000100110", --   94 -  376
      "00000010100101001011000000100110", --   95 -  380
      "00000000011001110100100000000110", --   96 -  384
      "00000010001101011011100000000110", --   97 -  388
      "00000000100001010101000000101011", --   98 -  392
      "00000010010100111100000000101011", --   99 -  396
      "00111100000010111011000100000110", --  100 -  400
      "00111100000110011011000100000110", --  101 -  404
      "00000000001000000110000000100111", --  102 -  408
      "00000001111000001101000000100111", --  103 -  412
      "00000000000000000000000000000000", --  104 -  416
      "00000000000000000000000000000000", --  105 -  420
      "00000000100010110110100000100001", --  106 -  424
      "00000010010110011101100000100001", --  107 -  428
      "00000000100000100111000000100100", --  108 -  432
      "00000010010100001110000000100100", --  109 -  436
      "00000001110010010011000000000111", --  110 -  440
      "00000011100101111010000000000111", --  111 -  444
      "00000000000010100000110101000011", --  112 -  448
      "00000000000110000111110101000011", --  113 -  452
      "00000001110010010001000000100110", --  114 -  456
      "00000011100101111000000000100110", --  115 -  460
      "00000001010011010100100000100001", --  116 -  464
      "00000011000110111011100000100001", --  117 -  468
      "00111100000010101111100001001000", --  118 -  472
      "00111100000110001111100001001000", --  119 -  476
      "00110000100011010010101000100001", --  120 -  480
      "00110010010110110010101000100001", --  121 -  484
      "00010101011110010000000100000001", --  122 -  488
      "10101100000010110000010000110100", --  123 -  492
      "00110000010010111110100101000110", --  124 -  496
      "00110010000110011110100101000110", --  125 -  500
      "00000000000001000010010101000011", --  126 -  504
      "00000000000100101001010101000011", --  127 -  508
      "10001100000000100000010000110100", --  128 -  512
      "10001100000100000000010000110100", --  129 -  516
      "00010100010100001111111111111110", --  130 -  520
      "00010101000101100000000011111000", --  131 -  524
      "10101100000010000000010000110100", --  132 -  528
      "00110000010010000000001011101110", --  133 -  532
      "00110010000101100000001011101110", --  134 -  536
      "00010100010100000000000011110100", --  135 -  540
      "10101100000000100000010000111000", --  136 -  544
      "00000000110001110001000000100011", --  137 -  548
      "00000010100101011000000000100011", --  138 -  552
      "00000000000000000000000000000000", --  139 -  556
      "00000000000000000000000000000000", --  140 -  560
      "00000000001000110011000000100010", --  141 -  564
      "00000001111100011010000000100010", --  142 -  568
      "00000001011000100011100000100101", --  143 -  572
      "00000011001100001010100000100101", --  144 -  576
      "00000001110010010000100000100111", --  145 -  580
      "00000011100101110111100000100111", --  146 -  584
      "00010100111101010000000011101000", --  147 -  588
      "10101100000001110000010000111100", --  148 -  592
      "00000000101011100011100000100101", --  149 -  596
      "00000010011111001010100000100101", --  150 -  600
      "10001100000001010000010000111100", --  151 -  604
      "10001100000100110000010000111100", --  152 -  608
      "00010100101100111111111111111110", --  153 -  612
      "00000000101000110111000000000110", --  154 -  616
      "00000010011100011110000000000110", --  155 -  620
      "00110001110000110110101000011011", --  156 -  624
      "00110011100100010110101000011011", --  157 -  628
      "00000001011000100111000000100101", --  158 -  632
      "00000011001100001110000000100101", --  159 -  636
      "00100000110010111011100111011001", --  160 -  640
      "00100010100110011011100111011001", --  161 -  644
      "00000000000010100001010101000011", --  162 -  648
      "00000000000110001000010101000011", --  163 -  652
      "00111100000001101011111011010101", --  164 -  656
      "00111100000101001011111011010101", --  165 -  660
      "10001100000010100000010000111000", --  166 -  664
      "10001100000110000000010000111000", --  167 -  668
      "00010101010110001111111111111110", --  168 -  672
      "00010100101100110000000011010010", --  169 -  676
      "10101100000001010000010000111000", --  170 -  680
      "00000001010001110010100000100101", --  171 -  684
      "00000011000101011001100000100101", --  172 -  688
      "00010100101100110000000011001110", --  173 -  692
      "10101100000001010000010000111100", --  174 -  696
      "00000000001000100010100000100000", --  175 -  700
      "00000001111100001001100000100000", --  176 -  704
      "00000000101011010000100000100001", --  177 -  708
      "00000010011110110111100000100001", --  178 -  712
      "00101100001000100110111101000101", --  179 -  716
      "00101101111100000110111101000101", --  180 -  720
      "00000001011000110010100000000111", --  181 -  724
      "00000011001100011001100000000111", --  182 -  728
      "00000001001001010110100000100100", --  183 -  732
      "00000010111100111101100000100100", --  184 -  736
      "00000000110000100000100000100101", --  185 -  740
      "00000010100100000111100000100101", --  186 -  744
      "00000001000000010001100000100110", --  187 -  748
      "00000010110011111000100000100110", --  188 -  752
      "00101101000010010011000111001011", --  189 -  756
      "00101110110101110011000111001011", --  190 -  760
      "10001100000001010000010000110100", --  191 -  764
      "10001100000100110000010000110100", --  192 -  768
      "00010100101100111111111111111110", --  193 -  772
      "00101000101001101100000010111011", --  194 -  776
      "00101010011101001100000010111011", --  195 -  780
      "00000000011010110001000000100001", --  196 -  784
      "00000010001110011000000000100001", --  197 -  788
      "00000000111011000000100000100110", --  198 -  792
      "00000010101110100111100000100110", --  199 -  796
      "00000000001011100100000000101011", --  200 -  800
      "00000001111111001011000000101011", --  201 -  804
      "00000000000000000000000000000000", --  202 -  808
      "00000000000000000000000000000000", --  203 -  812
      "00000001101001000101100000000111", --  204 -  816
      "00000011011100101100100000000111", --  205 -  820
      "00010100101100110000000010101101", --  206 -  824
      "10101100000001010000010000011100", --  207 -  828
      "00000001010010010011100000100110", --  208 -  832
      "00000011000101111010100000100110", --  209 -  836
      "00000000000000000000000000000000", --  210 -  840
      "00000000000000000000000000000000", --  211 -  844
      "00000000000001100110000111000010", --  212 -  848
      "00000000000101001101000111000010", --  213 -  852
      "00000000000000100000111001000011", --  214 -  856
      "00000000000100000111111001000011", --  215 -  860
      "00100101000011101001000110111000", --  216 -  864
      "00100110110111001001000110111000", --  217 -  868
      "10001100000001000000010000111000", --  218 -  872
      "10001100000100100000010000111000", --  219 -  876
      "00010100100100101111111111111110", --  220 -  880
      "00010100100100100000000010011110", --  221 -  884
      "10101100000001000000010000100000", --  222 -  888
      "00110100011011011111111000101001", --  223 -  892
      "00110110001110111111111000101001", --  224 -  896
      "00100001100001010010111110011100", --  225 -  900
      "00100011010100110010111110011100", --  226 -  904
      "10001100000010100000010000111100", --  227 -  908
      "10001100000110000000010000111100", --  228 -  912
      "00010101010110001111111111111110", --  229 -  916
      "00000001010011010100100000100001", --  230 -  920
      "00000011000110111011100000100001", --  231 -  924
      "00000000000000000000000000000000", --  232 -  928
      "00000000000000000000000000000000", --  233 -  932
      "00000001011000000011000000101011", --  234 -  936
      "00000011001000001010000000101011", --  235 -  940
      "00000001001000010001000000100101", --  236 -  944
      "00000010111011111000000000100101", --  237 -  948
      "00000000000000000000000000000000", --  238 -  952
      "00000000000000000000000000000000", --  239 -  956
      "00000001110000100100000000100111", --  240 -  960
      "00000011100100001011000000100111", --  241 -  964
      "00010100101100110000000010001001", --  242 -  968
      "10101100000001010000010000100100", --  243 -  972
      "00010100110101000000000010000111", --  244 -  976
      "10101100000001100000010000101000", --  245 -  980
      "00010100111101010000000010000101", --  246 -  984
      "10101100000001110000010000101100", --  247 -  988
      "00000000000000000000000000000000", --  248 -  992
      "00000000000000000000000000000000", --  249 -  996
      "00010101000101100000000010000001", --  250 - 1000
      "10101100000010000000010000110000", --  251 - 1004
      "00100011110111011111111100000110", --  252 - 1008
      "00010011101000000000000000010011", --  253 - 1012
      "00100011110111011111111000001100", --  254 - 1016
      "00010011101000000000000000010001", --  255 - 1020
      "00100011110111011111110100010010", --  256 - 1024
      "00010011101000000000000000001111", --  257 - 1028
      "00100011110111101111111111111111", --  258 - 1032
      "00100011111111111111111111111111", --  259 - 1036
      "00010111110111110000000001110111", --  260 - 1040
      "00011111111000001111111101001011", --  261 - 1044
      "00010000000000000000000100000010", --  262 - 1048
      "00000000000000000000000000000000", --  263 - 1052
      "00000000000000000000000000000000", --  264 - 1056
      "00000000000000000000000000000000", --  265 - 1060
      "00000000000000000000000000000000", --  266 - 1064
      "00000000000000000000000000000000", --  267 - 1068
      "00000000000000000000000000000000", --  268 - 1072
      "00000000000000000000000000000000", --  269 - 1076
      "00000000000000000000000000000000", --  270 - 1080
      "00000000000000000000000000000000", --  271 - 1084
      "10001100000111010000011110010100", --  272 - 1088
      "00011111101000000000000000000011", --  273 - 1092
      "00100000000111010000000000111100", --  274 - 1096
      "00010000000000000000000000000010", --  275 - 1100
      "00100000000111010000000000000000", --  276 - 1104
      "00010100001011110000000001100110", --  277 - 1108
      "10101111101000010000011100011100", --  278 - 1112
      "10001100000111010000011110010100", --  279 - 1116
      "00011111101000000000000000000011", --  280 - 1120
      "00100000000111010000000000111100", --  281 - 1124
      "00010000000000000000000000000010", --  282 - 1128
      "00100000000111010000000000000000", --  283 - 1132
      "00010100010100000000000001011111", --  284 - 1136
      "10101111101000100000011100100000", --  285 - 1140
      "10001100000111010000011110010100", --  286 - 1144
      "00011111101000000000000000000011", --  287 - 1148
      "00100000000111010000000000111100", --  288 - 1152
      "00010000000000000000000000000010", --  289 - 1156
      "00100000000111010000000000000000", --  290 - 1160
      "00010100011100010000000001011000", --  291 - 1164
      "10101111101000110000011100100100", --  292 - 1168
      "10001100000111010000011110010100", --  293 - 1172
      "00011111101000000000000000000011", --  294 - 1176
      "00100000000111010000000000111100", --  295 - 1180
      "00010000000000000000000000000010", --  296 - 1184
      "00100000000111010000000000000000", --  297 - 1188
      "00010100100100100000000001010001", --  298 - 1192
      "10101111101001000000011100101000", --  299 - 1196
      "10001100000111010000011110010100", --  300 - 1200
      "00011111101000000000000000000011", --  301 - 1204
      "00100000000111010000000000111100", --  302 - 1208
      "00010000000000000000000000000010", --  303 - 1212
      "00100000000111010000000000000000", --  304 - 1216
      "00010100101100110000000001001010", --  305 - 1220
      "10101111101001010000011100101100", --  306 - 1224
      "10001100000111010000011110010100", --  307 - 1228
      "00011111101000000000000000000011", --  308 - 1232
      "00100000000111010000000000111100", --  309 - 1236
      "00010000000000000000000000000010", --  310 - 1240
      "00100000000111010000000000000000", --  311 - 1244
      "00010100110101000000000001000011", --  312 - 1248
      "10101111101001100000011100110000", --  313 - 1252
      "10001100000111010000011110010100", --  314 - 1256
      "00011111101000000000000000000011", --  315 - 1260
      "00100000000111010000000000111100", --  316 - 1264
      "00010000000000000000000000000010", --  317 - 1268
      "00100000000111010000000000000000", --  318 - 1272
      "00010100111101010000000000111100", --  319 - 1276
      "10101111101001110000011100110100", --  320 - 1280
      "10001100000111010000011110010100", --  321 - 1284
      "00011111101000000000000000000011", --  322 - 1288
      "00100000000111010000000000111100", --  323 - 1292
      "00010000000000000000000000000010", --  324 - 1296
      "00100000000111010000000000000000", --  325 - 1300
      "00010101000101100000000000110101", --  326 - 1304
      "10101111101010000000011100111000", --  327 - 1308
      "10001100000111010000011110010100", --  328 - 1312
      "00011111101000000000000000000011", --  329 - 1316
      "00100000000111010000000000111100", --  330 - 1320
      "00010000000000000000000000000010", --  331 - 1324
      "00100000000111010000000000000000", --  332 - 1328
      "00010101001101110000000000101110", --  333 - 1332
      "10101111101010010000011100111100", --  334 - 1336
      "10001100000111010000011110010100", --  335 - 1340
      "00011111101000000000000000000011", --  336 - 1344
      "00100000000111010000000000111100", --  337 - 1348
      "00010000000000000000000000000010", --  338 - 1352
      "00100000000111010000000000000000", --  339 - 1356
      "00010101010110000000000000100111", --  340 - 1360
      "10101111101010100000011101000000", --  341 - 1364
      "10001100000111010000011110010100", --  342 - 1368
      "00011111101000000000000000000011", --  343 - 1372
      "00100000000111010000000000111100", --  344 - 1376
      "00010000000000000000000000000010", --  345 - 1380
      "00100000000111010000000000000000", --  346 - 1384
      "00010101011110010000000000100000", --  347 - 1388
      "10101111101010110000011101000100", --  348 - 1392
      "10001100000111010000011110010100", --  349 - 1396
      "00011111101000000000000000000011", --  350 - 1400
      "00100000000111010000000000111100", --  351 - 1404
      "00010000000000000000000000000010", --  352 - 1408
      "00100000000111010000000000000000", --  353 - 1412
      "00010101100110100000000000011001", --  354 - 1416
      "10101111101011000000011101001000", --  355 - 1420
      "10001100000111010000011110010100", --  356 - 1424
      "00011111101000000000000000000011", --  357 - 1428
      "00100000000111010000000000111100", --  358 - 1432
      "00010000000000000000000000000010", --  359 - 1436
      "00100000000111010000000000000000", --  360 - 1440
      "00010101101110110000000000010010", --  361 - 1444
      "10101111101011010000011101001100", --  362 - 1448
      "10001100000111010000011110010100", --  363 - 1452
      "00011111101000000000000000000011", --  364 - 1456
      "00100000000111010000000000111100", --  365 - 1460
      "00010000000000000000000000000010", --  366 - 1464
      "00100000000111010000000000000000", --  367 - 1468
      "00010101110111000000000000001011", --  368 - 1472
      "10101111101011100000011101010000", --  369 - 1476
      "10001100000111010000011110010100", --  370 - 1480
      "00011111101000000000000000000011", --  371 - 1484
      "00100000000111010000000000111100", --  372 - 1488
      "00010000000000000000000000000010", --  373 - 1492
      "00100000000111010000000000000000", --  374 - 1496
      "00010111110111110000000000000100", --  375 - 1500
      "10101111101111100000011101010100", --  376 - 1504
      "10101100000111010000011110010100", --  377 - 1508
      "00010000000000001111111110001000", --  378 - 1512
      "10001100000111010000011110010100", --  379 - 1516
      "10001111101000010000011100011100", --  380 - 1520
      "10001100000111010000011110010100", --  381 - 1524
      "10001111101011110000011100011100", --  382 - 1528
      "00010100001011111111111111111100", --  383 - 1532
      "10001100000111010000011110010100", --  384 - 1536
      "10001111101000100000011100100000", --  385 - 1540
      "10001100000111010000011110010100", --  386 - 1544
      "10001111101100000000011100100000", --  387 - 1548
      "00010100010100001111111111111100", --  388 - 1552
      "10001100000111010000011110010100", --  389 - 1556
      "10001111101000110000011100100100", --  390 - 1560
      "10001100000111010000011110010100", --  391 - 1564
      "10001111101100010000011100100100", --  392 - 1568
      "00010100011100011111111111111100", --  393 - 1572
      "10001100000111010000011110010100", --  394 - 1576
      "10001111101001000000011100101000", --  395 - 1580
      "10001100000111010000011110010100", --  396 - 1584
      "10001111101100100000011100101000", --  397 - 1588
      "00010100100100101111111111111100", --  398 - 1592
      "10001100000111010000011110010100", --  399 - 1596
      "10001111101001010000011100101100", --  400 - 1600
      "10001100000111010000011110010100", --  401 - 1604
      "10001111101100110000011100101100", --  402 - 1608
      "00010100101100111111111111111100", --  403 - 1612
      "10001100000111010000011110010100", --  404 - 1616
      "10001111101001100000011100110000", --  405 - 1620
      "10001100000111010000011110010100", --  406 - 1624
      "10001111101101000000011100110000", --  407 - 1628
      "00010100110101001111111111111100", --  408 - 1632
      "10001100000111010000011110010100", --  409 - 1636
      "10001111101001110000011100110100", --  410 - 1640
      "10001100000111010000011110010100", --  411 - 1644
      "10001111101101010000011100110100", --  412 - 1648
      "00010100111101011111111111111100", --  413 - 1652
      "10001100000111010000011110010100", --  414 - 1656
      "10001111101010000000011100111000", --  415 - 1660
      "10001100000111010000011110010100", --  416 - 1664
      "10001111101101100000011100111000", --  417 - 1668
      "00010101000101101111111111111100", --  418 - 1672
      "10001100000111010000011110010100", --  419 - 1676
      "10001111101010010000011100111100", --  420 - 1680
      "10001100000111010000011110010100", --  421 - 1684
      "10001111101101110000011100111100", --  422 - 1688
      "00010101001101111111111111111100", --  423 - 1692
      "10001100000111010000011110010100", --  424 - 1696
      "10001111101010100000011101000000", --  425 - 1700
      "10001100000111010000011110010100", --  426 - 1704
      "10001111101110000000011101000000", --  427 - 1708
      "00010101010110001111111111111100", --  428 - 1712
      "10001100000111010000011110010100", --  429 - 1716
      "10001111101010110000011101000100", --  430 - 1720
      "10001100000111010000011110010100", --  431 - 1724
      "10001111101110010000011101000100", --  432 - 1728
      "00010101011110011111111111111100", --  433 - 1732
      "10001100000111010000011110010100", --  434 - 1736
      "10001111101011000000011101001000", --  435 - 1740
      "10001100000111010000011110010100", --  436 - 1744
      "10001111101110100000011101001000", --  437 - 1748
      "00010101100110101111111111111100", --  438 - 1752
      "10001100000111010000011110010100", --  439 - 1756
      "10001111101011010000011101001100", --  440 - 1760
      "10001100000111010000011110010100", --  441 - 1764
      "10001111101110110000011101001100", --  442 - 1768
      "00010101101110111111111111111100", --  443 - 1772
      "10001100000111010000011110010100", --  444 - 1776
      "10001111101011100000011101010000", --  445 - 1780
      "10001100000111010000011110010100", --  446 - 1784
      "10001111101111000000011101010000", --  447 - 1788
      "00010101110111001111111111111100", --  448 - 1792
      "10001100000111010000011110010100", --  449 - 1796
      "10001111101111100000011101010100", --  450 - 1800
      "10001100000111010000011110010100", --  451 - 1804
      "10001111101111110000011101010100", --  452 - 1808
      "00010111110111111111111111111100", --  453 - 1812
      "00010000000000001111111100111100", --  454 - 1816
      "00000000000000000000000000000000", --  455 - 1820
      "00000000000000000000000000000000", --  456 - 1824
      "00000000000000000000000000000000", --  457 - 1828
      "00000000000000000000000000000000", --  458 - 1832
      "00000000000000000000000000000000", --  459 - 1836
      "00000000000000000000000000000000", --  460 - 1840
      "00000000000000000000000000000000", --  461 - 1844
      "00000000000000000000000000000000", --  462 - 1848
      "00000000000000000000000000000000", --  463 - 1852
      "00000000000000000000000000000000", --  464 - 1856
      "00000000000000000000000000000000", --  465 - 1860
      "00000000000000000000000000000000", --  466 - 1864
      "00000000000000000000000000000000", --  467 - 1868
      "00000000000000000000000000000000", --  468 - 1872
      "00000000000000000000000000000000", --  469 - 1876
      "00000000000000000000000000000000", --  470 - 1880
      "00000000000000000000000000000000", --  471 - 1884
      "00000000000000000000000000000000", --  472 - 1888
      "00000000000000000000000000000000", --  473 - 1892
      "00000000000000000000000000000000", --  474 - 1896
      "00000000000000000000000000000000", --  475 - 1900
      "00000000000000000000000000000000", --  476 - 1904
      "00000000000000000000000000000000", --  477 - 1908
      "00000000000000000000000000000000", --  478 - 1912
      "00000000000000000000000000000000", --  479 - 1916
      "00000000000000000000000000000000", --  480 - 1920
      "00000000000000000000000000000000", --  481 - 1924
      "00000000000000000000000000000000", --  482 - 1928
      "00000000000000000000000000000000", --  483 - 1932
      "00000000000000000000000000000000", --  484 - 1936
      "00000000000000000000001111100111", --  485 - 1940
      "00000000000000000000000000000000", --  486 - 1944
      "00000000000000000000000000000000", --  487 - 1948
      "00000000000000000000000000000000", --  488 - 1952
      "00000000000000000000000000000000", --  489 - 1956
      "00000000000000000000000000000000", --  490 - 1960
      "00000000000000000000000000000000", --  491 - 1964
      "00000000000000000000000000000000", --  492 - 1968
      "00000000000000000000000000000000", --  493 - 1972
      "00000000000000000000000000000000", --  494 - 1976
      "00000000000000000000000000000000", --  495 - 1980
      "00000000000000000000000000000000", --  496 - 1984
      "00000000000000000000000000000000", --  497 - 1988
      "00000000000000000000000000000000", --  498 - 1992
      "00000000000000000000000000000000", --  499 - 1996
      "00000000000000000000000000000000", --  500 - 2000
      "00000000000000000000000000000000", --  501 - 2004
      "00000000000000000000000000000000", --  502 - 2008
      "00000000000000000000000000000000", --  503 - 2012
      "00000000000000000000000000000000", --  504 - 2016
      "00000000000000000000000000000000", --  505 - 2020
      "00000000000000000000000000000000", --  506 - 2024
      "00000000000000000000000000000000", --  507 - 2028
      "00000000000000000000000000000000", --  508 - 2032
      "00000000000000000000000000000000", --  509 - 2036
      "00000000000000000000000000000000", --  510 - 2040
      "00000000000000000000000000000000", --  511 - 2044
      "00000000000000000000000000000000", --  512 - 2048
      "00000000000000000000000000000000", --  513 - 2052
      "00000000000000000000000000000000", --  514 - 2056
      "00000000000000000000000000000000", --  515 - 2060
      "00000000000000000000000000000000", --  516 - 2064
      "00000000000000000000000000000000", --  517 - 2068
      "00000000000000000000000000000000", --  518 - 2072
      "00000000000000000000000000000000", --  519 - 2076
      "00000000000000000000000000000000");--  520 - 2080

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000011110001011000110";
         f_reg(4) <= "00000000000000010001000000100011";
         f_reg(5) <= "00110000010000110010110010110100";
         f_reg(6) <= "00000000000000100010010111000011";
         f_reg(7) <= "00000000100000110010100000100101";
         f_reg(8) <= "00000000101001000011000000100111";
         f_reg(9) <= "00000000000001000011100000100000";
         f_reg(10) <= "00000000110001100100000000100110";
         f_reg(11) <= "00000000011001110100100000000110";
         f_reg(12) <= "00000000100001010101000000101011";
         f_reg(13) <= "00111100000010111011000100000110";
         f_reg(14) <= "00000000001000000110000000100111";
         f_reg(15) <= "00000000000000000000000000000000";
         f_reg(16) <= "00000000100010110110100000100001";
         f_reg(17) <= "00000000100000100111000000100100";
         f_reg(18) <= "00000001110010010111100000000111";
         f_reg(19) <= "00000000000010101000010101000011";
         f_reg(20) <= "00000001110010011000100000100110";
         f_reg(21) <= "00000001010011011001000000100001";
         f_reg(22) <= "00111100000100111111100001001000";
         f_reg(23) <= "00110000100101000010101000100001";
         f_reg(24) <= "00110010001101011110100101000110";
         f_reg(25) <= "00000000000001000010010101000011";
         f_reg(26) <= "00110001011101100000001011101110";
         f_reg(27) <= "00000001111001111011100000100011";
         f_reg(28) <= "00000000000000000000000000000000";
         f_reg(29) <= "00000010000000111100000000100010";
         f_reg(30) <= "00000010101101111100100000100101";
         f_reg(31) <= "00000001110100101101000000100111";
         f_reg(32) <= "00000000101011101101100000100101";
         f_reg(33) <= "00000011001000111110000000000110";
         f_reg(34) <= "00110011100111010110101000011011";
         f_reg(35) <= "00000010101101111111000000100101";
         f_reg(36) <= "00100011000001101011100111011001";
         f_reg(37) <= "00000000000100110000110101000011";
         f_reg(38) <= "00111100000000101011111011010101";
         f_reg(39) <= "00000001011110110100100000100101";
         f_reg(40) <= "00000011010000010101000000100000";
         f_reg(41) <= "00000001010101000110100000100001";
         f_reg(42) <= "00101101101100010110111101000101";
         f_reg(43) <= "00000000110111010111100000000111";
         f_reg(44) <= "00000010010011110011100000100100";
         f_reg(45) <= "00000000010100011000000000100101";
         f_reg(46) <= "00000010110100000010100000100110";
         f_reg(47) <= "00101110110011100011000111001011";
         f_reg(48) <= "00101001000000111100000010111011";
         f_reg(49) <= "00000000101001101110000000100001";
         f_reg(50) <= "00000011011011001010100000100110";
         f_reg(51) <= "00000010101111101011100000101011";
         f_reg(52) <= "00000000000000000000000000000000";
         f_reg(53) <= "00000000111001001100000000000111";
         f_reg(54) <= "10101100000010000000010000011100";
         f_reg(55) <= "00000001011011101001100000100110";
         f_reg(56) <= "00000000000000000000000000000000";
         f_reg(57) <= "00000000000000111101000111000010";
         f_reg(58) <= "00000000000111000000111001000011";
         f_reg(59) <= "00100110111010101001000110111000";
         f_reg(60) <= "10101100000110010000010000100000";
         f_reg(61) <= "00110100101101001111111000101001";
         f_reg(62) <= "00100011010011010010111110011100";
         f_reg(63) <= "00000001001101001110100000100001";
         f_reg(64) <= "00000000000000000000000000000000";
         f_reg(65) <= "00000011000000001001000000101011";
         f_reg(66) <= "00000011101000010111100000100101";
         f_reg(67) <= "00000000000000000000000000000000";
         f_reg(68) <= "00000001010011110001000000100111";
         f_reg(69) <= "10101100000011010000010000100100";
         f_reg(70) <= "10101100000100100000010000101000";
         f_reg(71) <= "10101100000100110000010000101100";
         f_reg(72) <= "00000000000000000000000000000000";
         f_reg(73) <= "10101100000000100000010000110000";
         f_reg(74) <= "00100011111111111111111111111111";
         f_reg(75) <= "00011111111000001111111110111000";
         f_reg(76) <= "00010000000000000000000110111101";
         f_reg(77) <= "00111100000111100000001111100111";
         f_reg(78) <= "00111100000111110000001111100111";
         f_reg(79) <= "00000000000111101111010000000010";
         f_reg(80) <= "00000000000111111111110000000010";
         f_reg(81) <= "00111100000000011110001011000110";
         f_reg(82) <= "00111100000011111110001011000110";
         f_reg(83) <= "00000000000000010001000000100011";
         f_reg(84) <= "00000000000011111000000000100011";
         f_reg(85) <= "00110000010000110010110010110100";
         f_reg(86) <= "00110010000100010010110010110100";
         f_reg(87) <= "00000000000000100010010111000011";
         f_reg(88) <= "00000000000100001001010111000011";
         f_reg(89) <= "00000000100000110010100000100101";
         f_reg(90) <= "00000010010100011001100000100101";
         f_reg(91) <= "00000000101001000011000000100111";
         f_reg(92) <= "00000010011100101010000000100111";
         f_reg(93) <= "00000000000001000011100000100000";
         f_reg(94) <= "00000000000100101010100000100000";
         f_reg(95) <= "00000000110001100100000000100110";
         f_reg(96) <= "00000010100101001011000000100110";
         f_reg(97) <= "00000000011001110100100000000110";
         f_reg(98) <= "00000010001101011011100000000110";
         f_reg(99) <= "00000000100001010101000000101011";
         f_reg(100) <= "00000010010100111100000000101011";
         f_reg(101) <= "00111100000010111011000100000110";
         f_reg(102) <= "00111100000110011011000100000110";
         f_reg(103) <= "00000000001000000110000000100111";
         f_reg(104) <= "00000001111000001101000000100111";
         f_reg(105) <= "00000000000000000000000000000000";
         f_reg(106) <= "00000000000000000000000000000000";
         f_reg(107) <= "00000000100010110110100000100001";
         f_reg(108) <= "00000010010110011101100000100001";
         f_reg(109) <= "00000000100000100111000000100100";
         f_reg(110) <= "00000010010100001110000000100100";
         f_reg(111) <= "00000001110010010011000000000111";
         f_reg(112) <= "00000011100101111010000000000111";
         f_reg(113) <= "00000000000010100000110101000011";
         f_reg(114) <= "00000000000110000111110101000011";
         f_reg(115) <= "00000001110010010001000000100110";
         f_reg(116) <= "00000011100101111000000000100110";
         f_reg(117) <= "00000001010011010100100000100001";
         f_reg(118) <= "00000011000110111011100000100001";
         f_reg(119) <= "00111100000010101111100001001000";
         f_reg(120) <= "00111100000110001111100001001000";
         f_reg(121) <= "00110000100011010010101000100001";
         f_reg(122) <= "00110010010110110010101000100001";
         f_reg(123) <= "00010101011110010000000100000001";
         f_reg(124) <= "10101100000010110000010000110100";
         f_reg(125) <= "00110000010010111110100101000110";
         f_reg(126) <= "00110010000110011110100101000110";
         f_reg(127) <= "00000000000001000010010101000011";
         f_reg(128) <= "00000000000100101001010101000011";
         f_reg(129) <= "10001100000000100000010000110100";
         f_reg(130) <= "10001100000100000000010000110100";
         f_reg(131) <= "00010100010100001111111111111110";
         f_reg(132) <= "00010101000101100000000011111000";
         f_reg(133) <= "10101100000010000000010000110100";
         f_reg(134) <= "00110000010010000000001011101110";
         f_reg(135) <= "00110010000101100000001011101110";
         f_reg(136) <= "00010100010100000000000011110100";
         f_reg(137) <= "10101100000000100000010000111000";
         f_reg(138) <= "00000000110001110001000000100011";
         f_reg(139) <= "00000010100101011000000000100011";
         f_reg(140) <= "00000000000000000000000000000000";
         f_reg(141) <= "00000000000000000000000000000000";
         f_reg(142) <= "00000000001000110011000000100010";
         f_reg(143) <= "00000001111100011010000000100010";
         f_reg(144) <= "00000001011000100011100000100101";
         f_reg(145) <= "00000011001100001010100000100101";
         f_reg(146) <= "00000001110010010000100000100111";
         f_reg(147) <= "00000011100101110111100000100111";
         f_reg(148) <= "00010100111101010000000011101000";
         f_reg(149) <= "10101100000001110000010000111100";
         f_reg(150) <= "00000000101011100011100000100101";
         f_reg(151) <= "00000010011111001010100000100101";
         f_reg(152) <= "10001100000001010000010000111100";
         f_reg(153) <= "10001100000100110000010000111100";
         f_reg(154) <= "00010100101100111111111111111110";
         f_reg(155) <= "00000000101000110111000000000110";
         f_reg(156) <= "00000010011100011110000000000110";
         f_reg(157) <= "00110001110000110110101000011011";
         f_reg(158) <= "00110011100100010110101000011011";
         f_reg(159) <= "00000001011000100111000000100101";
         f_reg(160) <= "00000011001100001110000000100101";
         f_reg(161) <= "00100000110010111011100111011001";
         f_reg(162) <= "00100010100110011011100111011001";
         f_reg(163) <= "00000000000010100001010101000011";
         f_reg(164) <= "00000000000110001000010101000011";
         f_reg(165) <= "00111100000001101011111011010101";
         f_reg(166) <= "00111100000101001011111011010101";
         f_reg(167) <= "10001100000010100000010000111000";
         f_reg(168) <= "10001100000110000000010000111000";
         f_reg(169) <= "00010101010110001111111111111110";
         f_reg(170) <= "00010100101100110000000011010010";
         f_reg(171) <= "10101100000001010000010000111000";
         f_reg(172) <= "00000001010001110010100000100101";
         f_reg(173) <= "00000011000101011001100000100101";
         f_reg(174) <= "00010100101100110000000011001110";
         f_reg(175) <= "10101100000001010000010000111100";
         f_reg(176) <= "00000000001000100010100000100000";
         f_reg(177) <= "00000001111100001001100000100000";
         f_reg(178) <= "00000000101011010000100000100001";
         f_reg(179) <= "00000010011110110111100000100001";
         f_reg(180) <= "00101100001000100110111101000101";
         f_reg(181) <= "00101101111100000110111101000101";
         f_reg(182) <= "00000001011000110010100000000111";
         f_reg(183) <= "00000011001100011001100000000111";
         f_reg(184) <= "00000001001001010110100000100100";
         f_reg(185) <= "00000010111100111101100000100100";
         f_reg(186) <= "00000000110000100000100000100101";
         f_reg(187) <= "00000010100100000111100000100101";
         f_reg(188) <= "00000001000000010001100000100110";
         f_reg(189) <= "00000010110011111000100000100110";
         f_reg(190) <= "00101101000010010011000111001011";
         f_reg(191) <= "00101110110101110011000111001011";
         f_reg(192) <= "10001100000001010000010000110100";
         f_reg(193) <= "10001100000100110000010000110100";
         f_reg(194) <= "00010100101100111111111111111110";
         f_reg(195) <= "00101000101001101100000010111011";
         f_reg(196) <= "00101010011101001100000010111011";
         f_reg(197) <= "00000000011010110001000000100001";
         f_reg(198) <= "00000010001110011000000000100001";
         f_reg(199) <= "00000000111011000000100000100110";
         f_reg(200) <= "00000010101110100111100000100110";
         f_reg(201) <= "00000000001011100100000000101011";
         f_reg(202) <= "00000001111111001011000000101011";
         f_reg(203) <= "00000000000000000000000000000000";
         f_reg(204) <= "00000000000000000000000000000000";
         f_reg(205) <= "00000001101001000101100000000111";
         f_reg(206) <= "00000011011100101100100000000111";
         f_reg(207) <= "00010100101100110000000010101101";
         f_reg(208) <= "10101100000001010000010000011100";
         f_reg(209) <= "00000001010010010011100000100110";
         f_reg(210) <= "00000011000101111010100000100110";
         f_reg(211) <= "00000000000000000000000000000000";
         f_reg(212) <= "00000000000000000000000000000000";
         f_reg(213) <= "00000000000001100110000111000010";
         f_reg(214) <= "00000000000101001101000111000010";
         f_reg(215) <= "00000000000000100000111001000011";
         f_reg(216) <= "00000000000100000111111001000011";
         f_reg(217) <= "00100101000011101001000110111000";
         f_reg(218) <= "00100110110111001001000110111000";
         f_reg(219) <= "10001100000001000000010000111000";
         f_reg(220) <= "10001100000100100000010000111000";
         f_reg(221) <= "00010100100100101111111111111110";
         f_reg(222) <= "00010100100100100000000010011110";
         f_reg(223) <= "10101100000001000000010000100000";
         f_reg(224) <= "00110100011011011111111000101001";
         f_reg(225) <= "00110110001110111111111000101001";
         f_reg(226) <= "00100001100001010010111110011100";
         f_reg(227) <= "00100011010100110010111110011100";
         f_reg(228) <= "10001100000010100000010000111100";
         f_reg(229) <= "10001100000110000000010000111100";
         f_reg(230) <= "00010101010110001111111111111110";
         f_reg(231) <= "00000001010011010100100000100001";
         f_reg(232) <= "00000011000110111011100000100001";
         f_reg(233) <= "00000000000000000000000000000000";
         f_reg(234) <= "00000000000000000000000000000000";
         f_reg(235) <= "00000001011000000011000000101011";
         f_reg(236) <= "00000011001000001010000000101011";
         f_reg(237) <= "00000001001000010001000000100101";
         f_reg(238) <= "00000010111011111000000000100101";
         f_reg(239) <= "00000000000000000000000000000000";
         f_reg(240) <= "00000000000000000000000000000000";
         f_reg(241) <= "00000001110000100100000000100111";
         f_reg(242) <= "00000011100100001011000000100111";
         f_reg(243) <= "00010100101100110000000010001001";
         f_reg(244) <= "10101100000001010000010000100100";
         f_reg(245) <= "00010100110101000000000010000111";
         f_reg(246) <= "10101100000001100000010000101000";
         f_reg(247) <= "00010100111101010000000010000101";
         f_reg(248) <= "10101100000001110000010000101100";
         f_reg(249) <= "00000000000000000000000000000000";
         f_reg(250) <= "00000000000000000000000000000000";
         f_reg(251) <= "00010101000101100000000010000001";
         f_reg(252) <= "10101100000010000000010000110000";
         f_reg(253) <= "00100011110111011111111100000110";
         f_reg(254) <= "00010011101000000000000000010011";
         f_reg(255) <= "00100011110111011111111000001100";
         f_reg(256) <= "00010011101000000000000000010001";
         f_reg(257) <= "00100011110111011111110100010010";
         f_reg(258) <= "00010011101000000000000000001111";
         f_reg(259) <= "00100011110111101111111111111111";
         f_reg(260) <= "00100011111111111111111111111111";
         f_reg(261) <= "00010111110111110000000001110111";
         f_reg(262) <= "00011111111000001111111101001011";
         f_reg(263) <= "00010000000000000000000100000010";
         f_reg(264) <= "00000000000000000000000000000000";
         f_reg(265) <= "00000000000000000000000000000000";
         f_reg(266) <= "00000000000000000000000000000000";
         f_reg(267) <= "00000000000000000000000000000000";
         f_reg(268) <= "00000000000000000000000000000000";
         f_reg(269) <= "00000000000000000000000000000000";
         f_reg(270) <= "00000000000000000000000000000000";
         f_reg(271) <= "00000000000000000000000000000000";
         f_reg(272) <= "00000000000000000000000000000000";
         f_reg(273) <= "10001100000111010000011110010100";
         f_reg(274) <= "00011111101000000000000000000011";
         f_reg(275) <= "00100000000111010000000000111100";
         f_reg(276) <= "00010000000000000000000000000010";
         f_reg(277) <= "00100000000111010000000000000000";
         f_reg(278) <= "00010100001011110000000001100110";
         f_reg(279) <= "10101111101000010000011100011100";
         f_reg(280) <= "10001100000111010000011110010100";
         f_reg(281) <= "00011111101000000000000000000011";
         f_reg(282) <= "00100000000111010000000000111100";
         f_reg(283) <= "00010000000000000000000000000010";
         f_reg(284) <= "00100000000111010000000000000000";
         f_reg(285) <= "00010100010100000000000001011111";
         f_reg(286) <= "10101111101000100000011100100000";
         f_reg(287) <= "10001100000111010000011110010100";
         f_reg(288) <= "00011111101000000000000000000011";
         f_reg(289) <= "00100000000111010000000000111100";
         f_reg(290) <= "00010000000000000000000000000010";
         f_reg(291) <= "00100000000111010000000000000000";
         f_reg(292) <= "00010100011100010000000001011000";
         f_reg(293) <= "10101111101000110000011100100100";
         f_reg(294) <= "10001100000111010000011110010100";
         f_reg(295) <= "00011111101000000000000000000011";
         f_reg(296) <= "00100000000111010000000000111100";
         f_reg(297) <= "00010000000000000000000000000010";
         f_reg(298) <= "00100000000111010000000000000000";
         f_reg(299) <= "00010100100100100000000001010001";
         f_reg(300) <= "10101111101001000000011100101000";
         f_reg(301) <= "10001100000111010000011110010100";
         f_reg(302) <= "00011111101000000000000000000011";
         f_reg(303) <= "00100000000111010000000000111100";
         f_reg(304) <= "00010000000000000000000000000010";
         f_reg(305) <= "00100000000111010000000000000000";
         f_reg(306) <= "00010100101100110000000001001010";
         f_reg(307) <= "10101111101001010000011100101100";
         f_reg(308) <= "10001100000111010000011110010100";
         f_reg(309) <= "00011111101000000000000000000011";
         f_reg(310) <= "00100000000111010000000000111100";
         f_reg(311) <= "00010000000000000000000000000010";
         f_reg(312) <= "00100000000111010000000000000000";
         f_reg(313) <= "00010100110101000000000001000011";
         f_reg(314) <= "10101111101001100000011100110000";
         f_reg(315) <= "10001100000111010000011110010100";
         f_reg(316) <= "00011111101000000000000000000011";
         f_reg(317) <= "00100000000111010000000000111100";
         f_reg(318) <= "00010000000000000000000000000010";
         f_reg(319) <= "00100000000111010000000000000000";
         f_reg(320) <= "00010100111101010000000000111100";
         f_reg(321) <= "10101111101001110000011100110100";
         f_reg(322) <= "10001100000111010000011110010100";
         f_reg(323) <= "00011111101000000000000000000011";
         f_reg(324) <= "00100000000111010000000000111100";
         f_reg(325) <= "00010000000000000000000000000010";
         f_reg(326) <= "00100000000111010000000000000000";
         f_reg(327) <= "00010101000101100000000000110101";
         f_reg(328) <= "10101111101010000000011100111000";
         f_reg(329) <= "10001100000111010000011110010100";
         f_reg(330) <= "00011111101000000000000000000011";
         f_reg(331) <= "00100000000111010000000000111100";
         f_reg(332) <= "00010000000000000000000000000010";
         f_reg(333) <= "00100000000111010000000000000000";
         f_reg(334) <= "00010101001101110000000000101110";
         f_reg(335) <= "10101111101010010000011100111100";
         f_reg(336) <= "10001100000111010000011110010100";
         f_reg(337) <= "00011111101000000000000000000011";
         f_reg(338) <= "00100000000111010000000000111100";
         f_reg(339) <= "00010000000000000000000000000010";
         f_reg(340) <= "00100000000111010000000000000000";
         f_reg(341) <= "00010101010110000000000000100111";
         f_reg(342) <= "10101111101010100000011101000000";
         f_reg(343) <= "10001100000111010000011110010100";
         f_reg(344) <= "00011111101000000000000000000011";
         f_reg(345) <= "00100000000111010000000000111100";
         f_reg(346) <= "00010000000000000000000000000010";
         f_reg(347) <= "00100000000111010000000000000000";
         f_reg(348) <= "00010101011110010000000000100000";
         f_reg(349) <= "10101111101010110000011101000100";
         f_reg(350) <= "10001100000111010000011110010100";
         f_reg(351) <= "00011111101000000000000000000011";
         f_reg(352) <= "00100000000111010000000000111100";
         f_reg(353) <= "00010000000000000000000000000010";
         f_reg(354) <= "00100000000111010000000000000000";
         f_reg(355) <= "00010101100110100000000000011001";
         f_reg(356) <= "10101111101011000000011101001000";
         f_reg(357) <= "10001100000111010000011110010100";
         f_reg(358) <= "00011111101000000000000000000011";
         f_reg(359) <= "00100000000111010000000000111100";
         f_reg(360) <= "00010000000000000000000000000010";
         f_reg(361) <= "00100000000111010000000000000000";
         f_reg(362) <= "00010101101110110000000000010010";
         f_reg(363) <= "10101111101011010000011101001100";
         f_reg(364) <= "10001100000111010000011110010100";
         f_reg(365) <= "00011111101000000000000000000011";
         f_reg(366) <= "00100000000111010000000000111100";
         f_reg(367) <= "00010000000000000000000000000010";
         f_reg(368) <= "00100000000111010000000000000000";
         f_reg(369) <= "00010101110111000000000000001011";
         f_reg(370) <= "10101111101011100000011101010000";
         f_reg(371) <= "10001100000111010000011110010100";
         f_reg(372) <= "00011111101000000000000000000011";
         f_reg(373) <= "00100000000111010000000000111100";
         f_reg(374) <= "00010000000000000000000000000010";
         f_reg(375) <= "00100000000111010000000000000000";
         f_reg(376) <= "00010111110111110000000000000100";
         f_reg(377) <= "10101111101111100000011101010100";
         f_reg(378) <= "10101100000111010000011110010100";
         f_reg(379) <= "00010000000000001111111110001000";
         f_reg(380) <= "10001100000111010000011110010100";
         f_reg(381) <= "10001111101000010000011100011100";
         f_reg(382) <= "10001100000111010000011110010100";
         f_reg(383) <= "10001111101011110000011100011100";
         f_reg(384) <= "00010100001011111111111111111100";
         f_reg(385) <= "10001100000111010000011110010100";
         f_reg(386) <= "10001111101000100000011100100000";
         f_reg(387) <= "10001100000111010000011110010100";
         f_reg(388) <= "10001111101100000000011100100000";
         f_reg(389) <= "00010100010100001111111111111100";
         f_reg(390) <= "10001100000111010000011110010100";
         f_reg(391) <= "10001111101000110000011100100100";
         f_reg(392) <= "10001100000111010000011110010100";
         f_reg(393) <= "10001111101100010000011100100100";
         f_reg(394) <= "00010100011100011111111111111100";
         f_reg(395) <= "10001100000111010000011110010100";
         f_reg(396) <= "10001111101001000000011100101000";
         f_reg(397) <= "10001100000111010000011110010100";
         f_reg(398) <= "10001111101100100000011100101000";
         f_reg(399) <= "00010100100100101111111111111100";
         f_reg(400) <= "10001100000111010000011110010100";
         f_reg(401) <= "10001111101001010000011100101100";
         f_reg(402) <= "10001100000111010000011110010100";
         f_reg(403) <= "10001111101100110000011100101100";
         f_reg(404) <= "00010100101100111111111111111100";
         f_reg(405) <= "10001100000111010000011110010100";
         f_reg(406) <= "10001111101001100000011100110000";
         f_reg(407) <= "10001100000111010000011110010100";
         f_reg(408) <= "10001111101101000000011100110000";
         f_reg(409) <= "00010100110101001111111111111100";
         f_reg(410) <= "10001100000111010000011110010100";
         f_reg(411) <= "10001111101001110000011100110100";
         f_reg(412) <= "10001100000111010000011110010100";
         f_reg(413) <= "10001111101101010000011100110100";
         f_reg(414) <= "00010100111101011111111111111100";
         f_reg(415) <= "10001100000111010000011110010100";
         f_reg(416) <= "10001111101010000000011100111000";
         f_reg(417) <= "10001100000111010000011110010100";
         f_reg(418) <= "10001111101101100000011100111000";
         f_reg(419) <= "00010101000101101111111111111100";
         f_reg(420) <= "10001100000111010000011110010100";
         f_reg(421) <= "10001111101010010000011100111100";
         f_reg(422) <= "10001100000111010000011110010100";
         f_reg(423) <= "10001111101101110000011100111100";
         f_reg(424) <= "00010101001101111111111111111100";
         f_reg(425) <= "10001100000111010000011110010100";
         f_reg(426) <= "10001111101010100000011101000000";
         f_reg(427) <= "10001100000111010000011110010100";
         f_reg(428) <= "10001111101110000000011101000000";
         f_reg(429) <= "00010101010110001111111111111100";
         f_reg(430) <= "10001100000111010000011110010100";
         f_reg(431) <= "10001111101010110000011101000100";
         f_reg(432) <= "10001100000111010000011110010100";
         f_reg(433) <= "10001111101110010000011101000100";
         f_reg(434) <= "00010101011110011111111111111100";
         f_reg(435) <= "10001100000111010000011110010100";
         f_reg(436) <= "10001111101011000000011101001000";
         f_reg(437) <= "10001100000111010000011110010100";
         f_reg(438) <= "10001111101110100000011101001000";
         f_reg(439) <= "00010101100110101111111111111100";
         f_reg(440) <= "10001100000111010000011110010100";
         f_reg(441) <= "10001111101011010000011101001100";
         f_reg(442) <= "10001100000111010000011110010100";
         f_reg(443) <= "10001111101110110000011101001100";
         f_reg(444) <= "00010101101110111111111111111100";
         f_reg(445) <= "10001100000111010000011110010100";
         f_reg(446) <= "10001111101011100000011101010000";
         f_reg(447) <= "10001100000111010000011110010100";
         f_reg(448) <= "10001111101111000000011101010000";
         f_reg(449) <= "00010101110111001111111111111100";
         f_reg(450) <= "10001100000111010000011110010100";
         f_reg(451) <= "10001111101111100000011101010100";
         f_reg(452) <= "10001100000111010000011110010100";
         f_reg(453) <= "10001111101111110000011101010100";
         f_reg(454) <= "00010111110111111111111111111100";
         f_reg(455) <= "00010000000000001111111100111100";
         f_reg(456) <= "00000000000000000000000000000000";
         f_reg(457) <= "00000000000000000000000000000000";
         f_reg(458) <= "00000000000000000000000000000000";
         f_reg(459) <= "00000000000000000000000000000000";
         f_reg(460) <= "00000000000000000000000000000000";
         f_reg(461) <= "00000000000000000000000000000000";
         f_reg(462) <= "00000000000000000000000000000000";
         f_reg(463) <= "00000000000000000000000000000000";
         f_reg(464) <= "00000000000000000000000000000000";
         f_reg(465) <= "00000000000000000000000000000000";
         f_reg(466) <= "00000000000000000000000000000000";
         f_reg(467) <= "00000000000000000000000000000000";
         f_reg(468) <= "00000000000000000000000000000000";
         f_reg(469) <= "00000000000000000000000000000000";
         f_reg(470) <= "00000000000000000000000000000000";
         f_reg(471) <= "00000000000000000000000000000000";
         f_reg(472) <= "00000000000000000000000000000000";
         f_reg(473) <= "00000000000000000000000000000000";
         f_reg(474) <= "00000000000000000000000000000000";
         f_reg(475) <= "00000000000000000000000000000000";
         f_reg(476) <= "00000000000000000000000000000000";
         f_reg(477) <= "00000000000000000000000000000000";
         f_reg(478) <= "00000000000000000000000000000000";
         f_reg(479) <= "00000000000000000000000000000000";
         f_reg(480) <= "00000000000000000000000000000000";
         f_reg(481) <= "00000000000000000000000000000000";
         f_reg(482) <= "00000000000000000000000000000000";
         f_reg(483) <= "00000000000000000000000000000000";
         f_reg(484) <= "00000000000000000000000000000000";
         f_reg(485) <= "00000000000000000000000000000000";
         f_reg(486) <= "00000000000000000000001111100111";
         f_reg(487) <= "00000000000000000000000000000000";
         f_reg(488) <= "00000000000000000000000000000000";
         f_reg(489) <= "00000000000000000000000000000000";
         f_reg(490) <= "00000000000000000000000000000000";
         f_reg(491) <= "00000000000000000000000000000000";
         f_reg(492) <= "00000000000000000000000000000000";
         f_reg(493) <= "00000000000000000000000000000000";
         f_reg(494) <= "00000000000000000000000000000000";
         f_reg(495) <= "00000000000000000000000000000000";
         f_reg(496) <= "00000000000000000000000000000000";
         f_reg(497) <= "00000000000000000000000000000000";
         f_reg(498) <= "00000000000000000000000000000000";
         f_reg(499) <= "00000000000000000000000000000000";
         f_reg(500) <= "00000000000000000000000000000000";
         f_reg(501) <= "00000000000000000000000000000000";
         f_reg(502) <= "00000000000000000000000000000000";
         f_reg(503) <= "00000000000000000000000000000000";
         f_reg(504) <= "00000000000000000000000000000000";
         f_reg(505) <= "00000000000000000000000000000000";
         f_reg(506) <= "00000000000000000000000000000000";
         f_reg(507) <= "00000000000000000000000000000000";
         f_reg(508) <= "00000000000000000000000000000000";
         f_reg(509) <= "00000000000000000000000000000000";
         f_reg(510) <= "00000000000000000000000000000000";
         f_reg(511) <= "00000000000000000000000000000000";
         f_reg(512) <= "00000000000000000000000000000000";
         f_reg(513) <= "00000000000000000000000000000000";
         f_reg(514) <= "00000000000000000000000000000000";
         f_reg(515) <= "00000000000000000000000000000000";
         f_reg(516) <= "00000000000000000000000000000000";
         f_reg(517) <= "00000000000000000000000000000000";
         f_reg(518) <= "00000000000000000000000000000000";
         f_reg(519) <= "00000000000000000000000000000000";
         f_reg(520) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 -7482
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SUBU R2 R0 R1
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- ANDI R3 R2 11444
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SRA R4 R2 23
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- OR R5 R4 R3
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- NOR R6 R5 R4
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- ADD R7 R0 R4
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- XOR R8 R6 R6
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- SRLV R9 R7 R3
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- SLTU R10 R4 R5
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- LUI R11 -20218
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- NOR R12 R1 R0
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- NOP
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- ADDU R13 R4 R11
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- AND R14 R4 R2
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- SRAV R15 R9 R14
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SRA R16 R10 21
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- XOR R17 R14 R9
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- ADDU R18 R10 R13
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- LUI R19 -1976
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- ANDI R20 R4 10785
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- ANDI R21 R17 -5818
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- SRA R4 R4 21
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- ANDI R22 R11 750
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- SUBU R23 R15 R7
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- NOP
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- SUB R24 R16 R3
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- OR R25 R21 R23
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- NOR R26 R14 R18
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- OR R27 R5 R14
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- SRLV R28 R3 R25
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- ANDI R29 R28 27163
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- OR R30 R21 R23
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- ADDI R6 R24 -17959
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- SRA R1 R19 21
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- LUI R2 -16683
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- OR R9 R11 R27
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- ADD R10 R26 R1
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- ADDU R13 R10 R20
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- SLTIU R17 R13 28485
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SRAV R15 R29 R6
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- AND R7 R18 R15
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- OR R16 R2 R17
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- XOR R5 R22 R16
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- SLTIU R14 R22 12747
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- SLTI R3 R8 -16197
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- ADDU R28 R5 R6
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- XOR R21 R27 R12
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SLTU R23 R21 R30
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- NOP
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- SRAV R24 R4 R7
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SW R8 R0 1052
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- XOR R19 R11 R14
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- NOP
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SRL R26 R3 7
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- SRA R1 R28 25
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- ADDIU R10 R23 -28232
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SW R25 R0 1056
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- ORI R20 R5 -471
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- ADDI R13 R26 12188
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- ADDU R29 R9 R20
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- NOP
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- SLTU R18 R24 R0
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- OR R15 R29 R1
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- NOP
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- NOR R2 R10 R15
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- SW R13 R0 1060
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SW R18 R0 1064
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- SW R19 R0 1068
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- NOP
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SW R2 R0 1072
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- BGTZ R31 -72
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- BEQ R0 R0 445
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- LUI R30 999
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- LUI R31 999
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- LUI R1 -7482
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- LUI R15 -7482
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SUBU R2 R0 R1
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- SUBU R16 R0 R15
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- ANDI R3 R2 11444
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- ANDI R17 R16 11444
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SRA R4 R2 23
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- SRA R18 R16 23
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- OR R5 R4 R3
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- OR R19 R18 R17
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- NOR R6 R5 R4
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- NOR R20 R19 R18
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- ADD R7 R0 R4
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- ADD R21 R0 R18
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- XOR R8 R6 R6
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- XOR R22 R20 R20
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SRLV R9 R7 R3
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SRLV R23 R21 R17
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- SLTU R10 R4 R5
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- SLTU R24 R18 R19
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- LUI R11 -20218
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- LUI R25 -20218
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- NOR R12 R1 R0
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- NOR R26 R15 R0
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- NOP
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- NOP
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- ADDU R13 R4 R11
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- ADDU R27 R18 R25
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- AND R14 R4 R2
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- AND R28 R18 R16
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- SRAV R6 R9 R14
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- SRAV R20 R23 R28
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- SRA R1 R10 21
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- SRA R15 R24 21
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- XOR R2 R14 R9
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- XOR R16 R28 R23
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- ADDU R9 R10 R13
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- ADDU R23 R24 R27
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- LUI R10 -1976
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- LUI R24 -1976
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- ANDI R13 R4 10785
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- ANDI R27 R18 10785
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- BNE R11 R25 257
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SW R11 R0 1076
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- ANDI R11 R2 -5818
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- ANDI R25 R16 -5818
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- SRA R4 R4 21
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SRA R18 R18 21
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- LW R2 R0 1076
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- LW R16 R0 1076
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- BNE R2 R16 -2
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- BNE R8 R22 248
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- SW R8 R0 1076
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- ANDI R8 R2 750
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- ANDI R22 R16 750
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- BNE R2 R16 244
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- SW R2 R0 1080
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SUBU R2 R6 R7
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- SUBU R16 R20 R21
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- NOP
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- NOP
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- SUB R6 R1 R3
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- SUB R20 R15 R17
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- OR R7 R11 R2
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- OR R21 R25 R16
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- NOR R1 R14 R9
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- NOR R15 R28 R23
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- BNE R7 R21 232
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- SW R7 R0 1084
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- OR R7 R5 R14
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- OR R21 R19 R28
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- LW R5 R0 1084
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- LW R19 R0 1084
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- BNE R5 R19 -2
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- SRLV R14 R3 R5
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- SRLV R28 R17 R19
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- ANDI R3 R14 27163
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- ANDI R17 R28 27163
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- OR R14 R11 R2
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- OR R28 R25 R16
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- ADDI R11 R6 -17959
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- ADDI R25 R20 -17959
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- SRA R2 R10 21
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- SRA R16 R24 21
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- LUI R6 -16683
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- LUI R20 -16683
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- LW R10 R0 1080
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- LW R24 R0 1080
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- BNE R10 R24 -2
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- BNE R5 R19 210
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- SW R5 R0 1080
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- OR R5 R10 R7
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- OR R19 R24 R21
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- BNE R5 R19 206
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- SW R5 R0 1084
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- ADD R5 R1 R2
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- ADD R19 R15 R16
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- ADDU R1 R5 R13
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- ADDU R15 R19 R27
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- SLTIU R2 R1 28485
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- SLTIU R16 R15 28485
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SRAV R5 R3 R11
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- SRAV R19 R17 R25
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- AND R13 R9 R5
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- AND R27 R23 R19
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- OR R1 R6 R2
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- OR R15 R20 R16
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- XOR R3 R8 R1
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- XOR R17 R22 R15
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- SLTIU R9 R8 12747
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- SLTIU R23 R22 12747
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- LW R5 R0 1076
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- LW R19 R0 1076
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- BNE R5 R19 -2
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- SLTI R6 R5 -16197
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- SLTI R20 R19 -16197
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- ADDU R2 R3 R11
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- ADDU R16 R17 R25
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- XOR R1 R7 R12
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- XOR R15 R21 R26
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- SLTU R8 R1 R14
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- SLTU R22 R15 R28
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- NOP
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- NOP
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- SRAV R11 R4 R13
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- SRAV R25 R18 R27
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- BNE R5 R19 173
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- SW R5 R0 1052
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- XOR R7 R10 R9
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- XOR R21 R24 R23
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- NOP
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- NOP
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- SRL R12 R6 7
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- SRL R26 R20 7
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- SRA R1 R2 25
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- SRA R15 R16 25
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- ADDIU R14 R8 -28232
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- ADDIU R28 R22 -28232
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- LW R4 R0 1080
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- LW R18 R0 1080
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- BNE R4 R18 -2
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- BNE R4 R18 158
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- SW R4 R0 1056
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- ORI R13 R3 -471
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- ORI R27 R17 -471
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- ADDI R5 R12 12188
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- ADDI R19 R26 12188
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- LW R10 R0 1084
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- LW R24 R0 1084
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- BNE R10 R24 -2
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- ADDU R9 R10 R13
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- ADDU R23 R24 R27
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- NOP
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- NOP
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- SLTU R6 R11 R0
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- SLTU R20 R25 R0
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- OR R2 R9 R1
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- OR R16 R23 R15
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- NOP
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- NOP
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- NOR R8 R14 R2
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- NOR R22 R28 R16
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- BNE R5 R19 137
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- SW R5 R0 1060
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- BNE R6 R20 135
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- SW R6 R0 1064
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- BNE R7 R21 133
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- SW R7 R0 1068
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- NOP
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- NOP
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- BNE R8 R22 129
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- SW R8 R0 1072
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- BEQ R29 R0 19
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- BEQ R29 R0 17
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- BEQ R29 R0 15
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- BNE R30 R31 119
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- BGTZ R31 -181
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- BEQ R0 R0 258
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- NOP
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- NOP
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- NOP
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- NOP
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- NOP
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- NOP
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- NOP
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- NOP
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- NOP
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- SW R1 R29 1820
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- SW R2 R29 1824
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- SW R3 R29 1828
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- SW R4 R29 1832
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- SW R5 R29 1836
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- SW R6 R29 1840
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- SW R7 R29 1844
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- SW R8 R29 1848
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- SW R9 R29 1852
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- SW R10 R29 1856
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- SW R11 R29 1860
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- SW R12 R29 1864
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- SW R13 R29 1868
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- SW R14 R29 1872
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- SW R30 R29 1876
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- SW R29 R0 1940
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- BEQ R0 R0 -120
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- LW R1 R29 1820
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- LW R15 R29 1820
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- LW R2 R29 1824
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- LW R16 R29 1824
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- LW R3 R29 1828
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- LW R17 R29 1828
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- LW R4 R29 1832
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- LW R18 R29 1832
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- LW R5 R29 1836
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- LW R19 R29 1836
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- LW R6 R29 1840
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- LW R20 R29 1840
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- LW R7 R29 1844
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- LW R21 R29 1844
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- LW R8 R29 1848
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- LW R22 R29 1848
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- LW R9 R29 1852
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- LW R23 R29 1852
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R10 R29 1856
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- LW R24 R29 1856
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- LW R11 R29 1860
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- LW R25 R29 1860
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- LW R12 R29 1864
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- LW R26 R29 1864
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- LW R13 R29 1868
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- LW R27 R29 1868
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- LW R14 R29 1872
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- LW R28 R29 1872
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- LW R30 R29 1876
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- LW R29 R0 1940
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- LW R31 R29 1876
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- BEQ R0 R0 -196
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- NOP
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- NOP
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- NOP
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- NOP
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- NOP
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- NOP
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- NOP
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- NOP
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- NOP
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- NOP
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- NOP
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- NOP
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- NOP
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- NOP
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- NOP
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- NOP
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- NOP
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- NOP
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- NOP
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- NOP
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- NOP
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- NOP
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- NOP
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- NOP
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- NOP
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- NOP
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- NOP
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- NOP
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- NOP
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- NOP
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- NOP
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- NOP
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- NOP
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- NOP
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- NOP
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- NOP
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- NOP
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- NOP
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- NOP
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- NOP
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- NOP
                        f_data <= f_reg(496);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(497) =>
                        -- NOP
                        f_data <= f_reg(497);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(498) =>
                        -- NOP
                        f_data <= f_reg(498);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(499) =>
                        -- NOP
                        f_data <= f_reg(499);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(500) =>
                        -- NOP
                        f_data <= f_reg(500);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(501) =>
                        -- NOP
                        f_data <= f_reg(501);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(502) =>
                        -- NOP
                        f_data <= f_reg(502);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(503) =>
                        -- NOP
                        f_data <= f_reg(503);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(504) =>
                        -- NOP
                        f_data <= f_reg(504);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(505) =>
                        -- NOP
                        f_data <= f_reg(505);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(506) =>
                        -- NOP
                        f_data <= f_reg(506);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(507) =>
                        -- NOP
                        f_data <= f_reg(507);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(508) =>
                        -- NOP
                        f_data <= f_reg(508);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(509) =>
                        -- NOP
                        f_data <= f_reg(509);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(510) =>
                        -- NOP
                        f_data <= f_reg(510);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(511) =>
                        -- NOP
                        f_data <= f_reg(511);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(512) =>
                        -- NOP
                        f_data <= f_reg(512);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(513) =>
                        -- NOP
                        f_data <= f_reg(513);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(514) =>
                        -- NOP
                        f_data <= f_reg(514);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(515) =>
                        -- NOP
                        f_data <= f_reg(515);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(516) =>
                        -- NOP
                        f_data <= f_reg(516);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(517) =>
                        -- NOP
                        f_data <= f_reg(517);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(518) =>
                        -- NOP
                        f_data <= f_reg(518);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(519) =>
                        -- NOP
                        f_data <= f_reg(519);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(520) =>
                        -- NOP
                        f_data <= f_reg(520);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(521) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011110001011000110";
                        f_reg(4) <= "00000000000000010001000000100011";
                        f_reg(5) <= "00110000010000110010110010110100";
                        f_reg(6) <= "00000000000000100010010111000011";
                        f_reg(7) <= "00000000100000110010100000100101";
                        f_reg(8) <= "00000000101001000011000000100111";
                        f_reg(9) <= "00000000000001000011100000100000";
                        f_reg(10) <= "00000000110001100100000000100110";
                        f_reg(11) <= "00000000011001110100100000000110";
                        f_reg(12) <= "00000000100001010101000000101011";
                        f_reg(13) <= "00111100000010111011000100000110";
                        f_reg(14) <= "00000000001000000110000000100111";
                        f_reg(15) <= "00000000000000000000000000000000";
                        f_reg(16) <= "00000000100010110110100000100001";
                        f_reg(17) <= "00000000100000100111000000100100";
                        f_reg(18) <= "00000001110010010111100000000111";
                        f_reg(19) <= "00000000000010101000010101000011";
                        f_reg(20) <= "00000001110010011000100000100110";
                        f_reg(21) <= "00000001010011011001000000100001";
                        f_reg(22) <= "00111100000100111111100001001000";
                        f_reg(23) <= "00110000100101000010101000100001";
                        f_reg(24) <= "00110010001101011110100101000110";
                        f_reg(25) <= "00000000000001000010010101000011";
                        f_reg(26) <= "00110001011101100000001011101110";
                        f_reg(27) <= "00000001111001111011100000100011";
                        f_reg(28) <= "00000000000000000000000000000000";
                        f_reg(29) <= "00000010000000111100000000100010";
                        f_reg(30) <= "00000010101101111100100000100101";
                        f_reg(31) <= "00000001110100101101000000100111";
                        f_reg(32) <= "00000000101011101101100000100101";
                        f_reg(33) <= "00000011001000111110000000000110";
                        f_reg(34) <= "00110011100111010110101000011011";
                        f_reg(35) <= "00000010101101111111000000100101";
                        f_reg(36) <= "00100011000001101011100111011001";
                        f_reg(37) <= "00000000000100110000110101000011";
                        f_reg(38) <= "00111100000000101011111011010101";
                        f_reg(39) <= "00000001011110110100100000100101";
                        f_reg(40) <= "00000011010000010101000000100000";
                        f_reg(41) <= "00000001010101000110100000100001";
                        f_reg(42) <= "00101101101100010110111101000101";
                        f_reg(43) <= "00000000110111010111100000000111";
                        f_reg(44) <= "00000010010011110011100000100100";
                        f_reg(45) <= "00000000010100011000000000100101";
                        f_reg(46) <= "00000010110100000010100000100110";
                        f_reg(47) <= "00101110110011100011000111001011";
                        f_reg(48) <= "00101001000000111100000010111011";
                        f_reg(49) <= "00000000101001101110000000100001";
                        f_reg(50) <= "00000011011011001010100000100110";
                        f_reg(51) <= "00000010101111101011100000101011";
                        f_reg(52) <= "00000000000000000000000000000000";
                        f_reg(53) <= "00000000111001001100000000000111";
                        f_reg(54) <= "10101100000010000000010000011100";
                        f_reg(55) <= "00000001011011101001100000100110";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000111101000111000010";
                        f_reg(58) <= "00000000000111000000111001000011";
                        f_reg(59) <= "00100110111010101001000110111000";
                        f_reg(60) <= "10101100000110010000010000100000";
                        f_reg(61) <= "00110100101101001111111000101001";
                        f_reg(62) <= "00100011010011010010111110011100";
                        f_reg(63) <= "00000001001101001110100000100001";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000011000000001001000000101011";
                        f_reg(66) <= "00000011101000010111100000100101";
                        f_reg(67) <= "00000000000000000000000000000000";
                        f_reg(68) <= "00000001010011110001000000100111";
                        f_reg(69) <= "10101100000011010000010000100100";
                        f_reg(70) <= "10101100000100100000010000101000";
                        f_reg(71) <= "10101100000100110000010000101100";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "10101100000000100000010000110000";
                        f_reg(74) <= "00100011111111111111111111111111";
                        f_reg(75) <= "00011111111000001111111110111000";
                        f_reg(76) <= "00010000000000000000000110111101";
                        f_reg(77) <= "00111100000111100000001111100111";
                        f_reg(78) <= "00111100000111110000001111100111";
                        f_reg(79) <= "00000000000111101111010000000010";
                        f_reg(80) <= "00000000000111111111110000000010";
                        f_reg(81) <= "00111100000000011110001011000110";
                        f_reg(82) <= "00111100000011111110001011000110";
                        f_reg(83) <= "00000000000000010001000000100011";
                        f_reg(84) <= "00000000000011111000000000100011";
                        f_reg(85) <= "00110000010000110010110010110100";
                        f_reg(86) <= "00110010000100010010110010110100";
                        f_reg(87) <= "00000000000000100010010111000011";
                        f_reg(88) <= "00000000000100001001010111000011";
                        f_reg(89) <= "00000000100000110010100000100101";
                        f_reg(90) <= "00000010010100011001100000100101";
                        f_reg(91) <= "00000000101001000011000000100111";
                        f_reg(92) <= "00000010011100101010000000100111";
                        f_reg(93) <= "00000000000001000011100000100000";
                        f_reg(94) <= "00000000000100101010100000100000";
                        f_reg(95) <= "00000000110001100100000000100110";
                        f_reg(96) <= "00000010100101001011000000100110";
                        f_reg(97) <= "00000000011001110100100000000110";
                        f_reg(98) <= "00000010001101011011100000000110";
                        f_reg(99) <= "00000000100001010101000000101011";
                        f_reg(100) <= "00000010010100111100000000101011";
                        f_reg(101) <= "00111100000010111011000100000110";
                        f_reg(102) <= "00111100000110011011000100000110";
                        f_reg(103) <= "00000000001000000110000000100111";
                        f_reg(104) <= "00000001111000001101000000100111";
                        f_reg(105) <= "00000000000000000000000000000000";
                        f_reg(106) <= "00000000000000000000000000000000";
                        f_reg(107) <= "00000000100010110110100000100001";
                        f_reg(108) <= "00000010010110011101100000100001";
                        f_reg(109) <= "00000000100000100111000000100100";
                        f_reg(110) <= "00000010010100001110000000100100";
                        f_reg(111) <= "00000001110010010011000000000111";
                        f_reg(112) <= "00000011100101111010000000000111";
                        f_reg(113) <= "00000000000010100000110101000011";
                        f_reg(114) <= "00000000000110000111110101000011";
                        f_reg(115) <= "00000001110010010001000000100110";
                        f_reg(116) <= "00000011100101111000000000100110";
                        f_reg(117) <= "00000001010011010100100000100001";
                        f_reg(118) <= "00000011000110111011100000100001";
                        f_reg(119) <= "00111100000010101111100001001000";
                        f_reg(120) <= "00111100000110001111100001001000";
                        f_reg(121) <= "00110000100011010010101000100001";
                        f_reg(122) <= "00110010010110110010101000100001";
                        f_reg(123) <= "00010101011110010000000100000001";
                        f_reg(124) <= "10101100000010110000010000110100";
                        f_reg(125) <= "00110000010010111110100101000110";
                        f_reg(126) <= "00110010000110011110100101000110";
                        f_reg(127) <= "00000000000001000010010101000011";
                        f_reg(128) <= "00000000000100101001010101000011";
                        f_reg(129) <= "10001100000000100000010000110100";
                        f_reg(130) <= "10001100000100000000010000110100";
                        f_reg(131) <= "00010100010100001111111111111110";
                        f_reg(132) <= "00010101000101100000000011111000";
                        f_reg(133) <= "10101100000010000000010000110100";
                        f_reg(134) <= "00110000010010000000001011101110";
                        f_reg(135) <= "00110010000101100000001011101110";
                        f_reg(136) <= "00010100010100000000000011110100";
                        f_reg(137) <= "10101100000000100000010000111000";
                        f_reg(138) <= "00000000110001110001000000100011";
                        f_reg(139) <= "00000010100101011000000000100011";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000000000000000000000000000";
                        f_reg(142) <= "00000000001000110011000000100010";
                        f_reg(143) <= "00000001111100011010000000100010";
                        f_reg(144) <= "00000001011000100011100000100101";
                        f_reg(145) <= "00000011001100001010100000100101";
                        f_reg(146) <= "00000001110010010000100000100111";
                        f_reg(147) <= "00000011100101110111100000100111";
                        f_reg(148) <= "00010100111101010000000011101000";
                        f_reg(149) <= "10101100000001110000010000111100";
                        f_reg(150) <= "00000000101011100011100000100101";
                        f_reg(151) <= "00000010011111001010100000100101";
                        f_reg(152) <= "10001100000001010000010000111100";
                        f_reg(153) <= "10001100000100110000010000111100";
                        f_reg(154) <= "00010100101100111111111111111110";
                        f_reg(155) <= "00000000101000110111000000000110";
                        f_reg(156) <= "00000010011100011110000000000110";
                        f_reg(157) <= "00110001110000110110101000011011";
                        f_reg(158) <= "00110011100100010110101000011011";
                        f_reg(159) <= "00000001011000100111000000100101";
                        f_reg(160) <= "00000011001100001110000000100101";
                        f_reg(161) <= "00100000110010111011100111011001";
                        f_reg(162) <= "00100010100110011011100111011001";
                        f_reg(163) <= "00000000000010100001010101000011";
                        f_reg(164) <= "00000000000110001000010101000011";
                        f_reg(165) <= "00111100000001101011111011010101";
                        f_reg(166) <= "00111100000101001011111011010101";
                        f_reg(167) <= "10001100000010100000010000111000";
                        f_reg(168) <= "10001100000110000000010000111000";
                        f_reg(169) <= "00010101010110001111111111111110";
                        f_reg(170) <= "00010100101100110000000011010010";
                        f_reg(171) <= "10101100000001010000010000111000";
                        f_reg(172) <= "00000001010001110010100000100101";
                        f_reg(173) <= "00000011000101011001100000100101";
                        f_reg(174) <= "00010100101100110000000011001110";
                        f_reg(175) <= "10101100000001010000010000111100";
                        f_reg(176) <= "00000000001000100010100000100000";
                        f_reg(177) <= "00000001111100001001100000100000";
                        f_reg(178) <= "00000000101011010000100000100001";
                        f_reg(179) <= "00000010011110110111100000100001";
                        f_reg(180) <= "00101100001000100110111101000101";
                        f_reg(181) <= "00101101111100000110111101000101";
                        f_reg(182) <= "00000001011000110010100000000111";
                        f_reg(183) <= "00000011001100011001100000000111";
                        f_reg(184) <= "00000001001001010110100000100100";
                        f_reg(185) <= "00000010111100111101100000100100";
                        f_reg(186) <= "00000000110000100000100000100101";
                        f_reg(187) <= "00000010100100000111100000100101";
                        f_reg(188) <= "00000001000000010001100000100110";
                        f_reg(189) <= "00000010110011111000100000100110";
                        f_reg(190) <= "00101101000010010011000111001011";
                        f_reg(191) <= "00101110110101110011000111001011";
                        f_reg(192) <= "10001100000001010000010000110100";
                        f_reg(193) <= "10001100000100110000010000110100";
                        f_reg(194) <= "00010100101100111111111111111110";
                        f_reg(195) <= "00101000101001101100000010111011";
                        f_reg(196) <= "00101010011101001100000010111011";
                        f_reg(197) <= "00000000011010110001000000100001";
                        f_reg(198) <= "00000010001110011000000000100001";
                        f_reg(199) <= "00000000111011000000100000100110";
                        f_reg(200) <= "00000010101110100111100000100110";
                        f_reg(201) <= "00000000001011100100000000101011";
                        f_reg(202) <= "00000001111111001011000000101011";
                        f_reg(203) <= "00000000000000000000000000000000";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000001101001000101100000000111";
                        f_reg(206) <= "00000011011100101100100000000111";
                        f_reg(207) <= "00010100101100110000000010101101";
                        f_reg(208) <= "10101100000001010000010000011100";
                        f_reg(209) <= "00000001010010010011100000100110";
                        f_reg(210) <= "00000011000101111010100000100110";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000001100110000111000010";
                        f_reg(214) <= "00000000000101001101000111000010";
                        f_reg(215) <= "00000000000000100000111001000011";
                        f_reg(216) <= "00000000000100000111111001000011";
                        f_reg(217) <= "00100101000011101001000110111000";
                        f_reg(218) <= "00100110110111001001000110111000";
                        f_reg(219) <= "10001100000001000000010000111000";
                        f_reg(220) <= "10001100000100100000010000111000";
                        f_reg(221) <= "00010100100100101111111111111110";
                        f_reg(222) <= "00010100100100100000000010011110";
                        f_reg(223) <= "10101100000001000000010000100000";
                        f_reg(224) <= "00110100011011011111111000101001";
                        f_reg(225) <= "00110110001110111111111000101001";
                        f_reg(226) <= "00100001100001010010111110011100";
                        f_reg(227) <= "00100011010100110010111110011100";
                        f_reg(228) <= "10001100000010100000010000111100";
                        f_reg(229) <= "10001100000110000000010000111100";
                        f_reg(230) <= "00010101010110001111111111111110";
                        f_reg(231) <= "00000001010011010100100000100001";
                        f_reg(232) <= "00000011000110111011100000100001";
                        f_reg(233) <= "00000000000000000000000000000000";
                        f_reg(234) <= "00000000000000000000000000000000";
                        f_reg(235) <= "00000001011000000011000000101011";
                        f_reg(236) <= "00000011001000001010000000101011";
                        f_reg(237) <= "00000001001000010001000000100101";
                        f_reg(238) <= "00000010111011111000000000100101";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000001110000100100000000100111";
                        f_reg(242) <= "00000011100100001011000000100111";
                        f_reg(243) <= "00010100101100110000000010001001";
                        f_reg(244) <= "10101100000001010000010000100100";
                        f_reg(245) <= "00010100110101000000000010000111";
                        f_reg(246) <= "10101100000001100000010000101000";
                        f_reg(247) <= "00010100111101010000000010000101";
                        f_reg(248) <= "10101100000001110000010000101100";
                        f_reg(249) <= "00000000000000000000000000000000";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00010101000101100000000010000001";
                        f_reg(252) <= "10101100000010000000010000110000";
                        f_reg(253) <= "00100011110111011111111100000110";
                        f_reg(254) <= "00010011101000000000000000010011";
                        f_reg(255) <= "00100011110111011111111000001100";
                        f_reg(256) <= "00010011101000000000000000010001";
                        f_reg(257) <= "00100011110111011111110100010010";
                        f_reg(258) <= "00010011101000000000000000001111";
                        f_reg(259) <= "00100011110111101111111111111111";
                        f_reg(260) <= "00100011111111111111111111111111";
                        f_reg(261) <= "00010111110111110000000001110111";
                        f_reg(262) <= "00011111111000001111111101001011";
                        f_reg(263) <= "00010000000000000000000100000010";
                        f_reg(264) <= "00000000000000000000000000000000";
                        f_reg(265) <= "00000000000000000000000000000000";
                        f_reg(266) <= "00000000000000000000000000000000";
                        f_reg(267) <= "00000000000000000000000000000000";
                        f_reg(268) <= "00000000000000000000000000000000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "10001100000111010000011110010100";
                        f_reg(274) <= "00011111101000000000000000000011";
                        f_reg(275) <= "00100000000111010000000000111100";
                        f_reg(276) <= "00010000000000000000000000000010";
                        f_reg(277) <= "00100000000111010000000000000000";
                        f_reg(278) <= "00010100001011110000000001100110";
                        f_reg(279) <= "10101111101000010000011100011100";
                        f_reg(280) <= "10001100000111010000011110010100";
                        f_reg(281) <= "00011111101000000000000000000011";
                        f_reg(282) <= "00100000000111010000000000111100";
                        f_reg(283) <= "00010000000000000000000000000010";
                        f_reg(284) <= "00100000000111010000000000000000";
                        f_reg(285) <= "00010100010100000000000001011111";
                        f_reg(286) <= "10101111101000100000011100100000";
                        f_reg(287) <= "10001100000111010000011110010100";
                        f_reg(288) <= "00011111101000000000000000000011";
                        f_reg(289) <= "00100000000111010000000000111100";
                        f_reg(290) <= "00010000000000000000000000000010";
                        f_reg(291) <= "00100000000111010000000000000000";
                        f_reg(292) <= "00010100011100010000000001011000";
                        f_reg(293) <= "10101111101000110000011100100100";
                        f_reg(294) <= "10001100000111010000011110010100";
                        f_reg(295) <= "00011111101000000000000000000011";
                        f_reg(296) <= "00100000000111010000000000111100";
                        f_reg(297) <= "00010000000000000000000000000010";
                        f_reg(298) <= "00100000000111010000000000000000";
                        f_reg(299) <= "00010100100100100000000001010001";
                        f_reg(300) <= "10101111101001000000011100101000";
                        f_reg(301) <= "10001100000111010000011110010100";
                        f_reg(302) <= "00011111101000000000000000000011";
                        f_reg(303) <= "00100000000111010000000000111100";
                        f_reg(304) <= "00010000000000000000000000000010";
                        f_reg(305) <= "00100000000111010000000000000000";
                        f_reg(306) <= "00010100101100110000000001001010";
                        f_reg(307) <= "10101111101001010000011100101100";
                        f_reg(308) <= "10001100000111010000011110010100";
                        f_reg(309) <= "00011111101000000000000000000011";
                        f_reg(310) <= "00100000000111010000000000111100";
                        f_reg(311) <= "00010000000000000000000000000010";
                        f_reg(312) <= "00100000000111010000000000000000";
                        f_reg(313) <= "00010100110101000000000001000011";
                        f_reg(314) <= "10101111101001100000011100110000";
                        f_reg(315) <= "10001100000111010000011110010100";
                        f_reg(316) <= "00011111101000000000000000000011";
                        f_reg(317) <= "00100000000111010000000000111100";
                        f_reg(318) <= "00010000000000000000000000000010";
                        f_reg(319) <= "00100000000111010000000000000000";
                        f_reg(320) <= "00010100111101010000000000111100";
                        f_reg(321) <= "10101111101001110000011100110100";
                        f_reg(322) <= "10001100000111010000011110010100";
                        f_reg(323) <= "00011111101000000000000000000011";
                        f_reg(324) <= "00100000000111010000000000111100";
                        f_reg(325) <= "00010000000000000000000000000010";
                        f_reg(326) <= "00100000000111010000000000000000";
                        f_reg(327) <= "00010101000101100000000000110101";
                        f_reg(328) <= "10101111101010000000011100111000";
                        f_reg(329) <= "10001100000111010000011110010100";
                        f_reg(330) <= "00011111101000000000000000000011";
                        f_reg(331) <= "00100000000111010000000000111100";
                        f_reg(332) <= "00010000000000000000000000000010";
                        f_reg(333) <= "00100000000111010000000000000000";
                        f_reg(334) <= "00010101001101110000000000101110";
                        f_reg(335) <= "10101111101010010000011100111100";
                        f_reg(336) <= "10001100000111010000011110010100";
                        f_reg(337) <= "00011111101000000000000000000011";
                        f_reg(338) <= "00100000000111010000000000111100";
                        f_reg(339) <= "00010000000000000000000000000010";
                        f_reg(340) <= "00100000000111010000000000000000";
                        f_reg(341) <= "00010101010110000000000000100111";
                        f_reg(342) <= "10101111101010100000011101000000";
                        f_reg(343) <= "10001100000111010000011110010100";
                        f_reg(344) <= "00011111101000000000000000000011";
                        f_reg(345) <= "00100000000111010000000000111100";
                        f_reg(346) <= "00010000000000000000000000000010";
                        f_reg(347) <= "00100000000111010000000000000000";
                        f_reg(348) <= "00010101011110010000000000100000";
                        f_reg(349) <= "10101111101010110000011101000100";
                        f_reg(350) <= "10001100000111010000011110010100";
                        f_reg(351) <= "00011111101000000000000000000011";
                        f_reg(352) <= "00100000000111010000000000111100";
                        f_reg(353) <= "00010000000000000000000000000010";
                        f_reg(354) <= "00100000000111010000000000000000";
                        f_reg(355) <= "00010101100110100000000000011001";
                        f_reg(356) <= "10101111101011000000011101001000";
                        f_reg(357) <= "10001100000111010000011110010100";
                        f_reg(358) <= "00011111101000000000000000000011";
                        f_reg(359) <= "00100000000111010000000000111100";
                        f_reg(360) <= "00010000000000000000000000000010";
                        f_reg(361) <= "00100000000111010000000000000000";
                        f_reg(362) <= "00010101101110110000000000010010";
                        f_reg(363) <= "10101111101011010000011101001100";
                        f_reg(364) <= "10001100000111010000011110010100";
                        f_reg(365) <= "00011111101000000000000000000011";
                        f_reg(366) <= "00100000000111010000000000111100";
                        f_reg(367) <= "00010000000000000000000000000010";
                        f_reg(368) <= "00100000000111010000000000000000";
                        f_reg(369) <= "00010101110111000000000000001011";
                        f_reg(370) <= "10101111101011100000011101010000";
                        f_reg(371) <= "10001100000111010000011110010100";
                        f_reg(372) <= "00011111101000000000000000000011";
                        f_reg(373) <= "00100000000111010000000000111100";
                        f_reg(374) <= "00010000000000000000000000000010";
                        f_reg(375) <= "00100000000111010000000000000000";
                        f_reg(376) <= "00010111110111110000000000000100";
                        f_reg(377) <= "10101111101111100000011101010100";
                        f_reg(378) <= "10101100000111010000011110010100";
                        f_reg(379) <= "00010000000000001111111110001000";
                        f_reg(380) <= "10001100000111010000011110010100";
                        f_reg(381) <= "10001111101000010000011100011100";
                        f_reg(382) <= "10001100000111010000011110010100";
                        f_reg(383) <= "10001111101011110000011100011100";
                        f_reg(384) <= "00010100001011111111111111111100";
                        f_reg(385) <= "10001100000111010000011110010100";
                        f_reg(386) <= "10001111101000100000011100100000";
                        f_reg(387) <= "10001100000111010000011110010100";
                        f_reg(388) <= "10001111101100000000011100100000";
                        f_reg(389) <= "00010100010100001111111111111100";
                        f_reg(390) <= "10001100000111010000011110010100";
                        f_reg(391) <= "10001111101000110000011100100100";
                        f_reg(392) <= "10001100000111010000011110010100";
                        f_reg(393) <= "10001111101100010000011100100100";
                        f_reg(394) <= "00010100011100011111111111111100";
                        f_reg(395) <= "10001100000111010000011110010100";
                        f_reg(396) <= "10001111101001000000011100101000";
                        f_reg(397) <= "10001100000111010000011110010100";
                        f_reg(398) <= "10001111101100100000011100101000";
                        f_reg(399) <= "00010100100100101111111111111100";
                        f_reg(400) <= "10001100000111010000011110010100";
                        f_reg(401) <= "10001111101001010000011100101100";
                        f_reg(402) <= "10001100000111010000011110010100";
                        f_reg(403) <= "10001111101100110000011100101100";
                        f_reg(404) <= "00010100101100111111111111111100";
                        f_reg(405) <= "10001100000111010000011110010100";
                        f_reg(406) <= "10001111101001100000011100110000";
                        f_reg(407) <= "10001100000111010000011110010100";
                        f_reg(408) <= "10001111101101000000011100110000";
                        f_reg(409) <= "00010100110101001111111111111100";
                        f_reg(410) <= "10001100000111010000011110010100";
                        f_reg(411) <= "10001111101001110000011100110100";
                        f_reg(412) <= "10001100000111010000011110010100";
                        f_reg(413) <= "10001111101101010000011100110100";
                        f_reg(414) <= "00010100111101011111111111111100";
                        f_reg(415) <= "10001100000111010000011110010100";
                        f_reg(416) <= "10001111101010000000011100111000";
                        f_reg(417) <= "10001100000111010000011110010100";
                        f_reg(418) <= "10001111101101100000011100111000";
                        f_reg(419) <= "00010101000101101111111111111100";
                        f_reg(420) <= "10001100000111010000011110010100";
                        f_reg(421) <= "10001111101010010000011100111100";
                        f_reg(422) <= "10001100000111010000011110010100";
                        f_reg(423) <= "10001111101101110000011100111100";
                        f_reg(424) <= "00010101001101111111111111111100";
                        f_reg(425) <= "10001100000111010000011110010100";
                        f_reg(426) <= "10001111101010100000011101000000";
                        f_reg(427) <= "10001100000111010000011110010100";
                        f_reg(428) <= "10001111101110000000011101000000";
                        f_reg(429) <= "00010101010110001111111111111100";
                        f_reg(430) <= "10001100000111010000011110010100";
                        f_reg(431) <= "10001111101010110000011101000100";
                        f_reg(432) <= "10001100000111010000011110010100";
                        f_reg(433) <= "10001111101110010000011101000100";
                        f_reg(434) <= "00010101011110011111111111111100";
                        f_reg(435) <= "10001100000111010000011110010100";
                        f_reg(436) <= "10001111101011000000011101001000";
                        f_reg(437) <= "10001100000111010000011110010100";
                        f_reg(438) <= "10001111101110100000011101001000";
                        f_reg(439) <= "00010101100110101111111111111100";
                        f_reg(440) <= "10001100000111010000011110010100";
                        f_reg(441) <= "10001111101011010000011101001100";
                        f_reg(442) <= "10001100000111010000011110010100";
                        f_reg(443) <= "10001111101110110000011101001100";
                        f_reg(444) <= "00010101101110111111111111111100";
                        f_reg(445) <= "10001100000111010000011110010100";
                        f_reg(446) <= "10001111101011100000011101010000";
                        f_reg(447) <= "10001100000111010000011110010100";
                        f_reg(448) <= "10001111101111000000011101010000";
                        f_reg(449) <= "00010101110111001111111111111100";
                        f_reg(450) <= "10001100000111010000011110010100";
                        f_reg(451) <= "10001111101111100000011101010100";
                        f_reg(452) <= "10001100000111010000011110010100";
                        f_reg(453) <= "10001111101111110000011101010100";
                        f_reg(454) <= "00010111110111111111111111111100";
                        f_reg(455) <= "00010000000000001111111100111100";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000001111100111";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011110001011000110";
                        f_reg(4) <= "00000000000000010001000000100011";
                        f_reg(5) <= "00110000010000110010110010110100";
                        f_reg(6) <= "00000000000000100010010111000011";
                        f_reg(7) <= "00000000100000110010100000100101";
                        f_reg(8) <= "00000000101001000011000000100111";
                        f_reg(9) <= "00000000000001000011100000100000";
                        f_reg(10) <= "00000000110001100100000000100110";
                        f_reg(11) <= "00000000011001110100100000000110";
                        f_reg(12) <= "00000000100001010101000000101011";
                        f_reg(13) <= "00111100000010111011000100000110";
                        f_reg(14) <= "00000000001000000110000000100111";
                        f_reg(15) <= "00000000000000000000000000000000";
                        f_reg(16) <= "00000000100010110110100000100001";
                        f_reg(17) <= "00000000100000100111000000100100";
                        f_reg(18) <= "00000001110010010111100000000111";
                        f_reg(19) <= "00000000000010101000010101000011";
                        f_reg(20) <= "00000001110010011000100000100110";
                        f_reg(21) <= "00000001010011011001000000100001";
                        f_reg(22) <= "00111100000100111111100001001000";
                        f_reg(23) <= "00110000100101000010101000100001";
                        f_reg(24) <= "00110010001101011110100101000110";
                        f_reg(25) <= "00000000000001000010010101000011";
                        f_reg(26) <= "00110001011101100000001011101110";
                        f_reg(27) <= "00000001111001111011100000100011";
                        f_reg(28) <= "00000000000000000000000000000000";
                        f_reg(29) <= "00000010000000111100000000100010";
                        f_reg(30) <= "00000010101101111100100000100101";
                        f_reg(31) <= "00000001110100101101000000100111";
                        f_reg(32) <= "00000000101011101101100000100101";
                        f_reg(33) <= "00000011001000111110000000000110";
                        f_reg(34) <= "00110011100111010110101000011011";
                        f_reg(35) <= "00000010101101111111000000100101";
                        f_reg(36) <= "00100011000001101011100111011001";
                        f_reg(37) <= "00000000000100110000110101000011";
                        f_reg(38) <= "00111100000000101011111011010101";
                        f_reg(39) <= "00000001011110110100100000100101";
                        f_reg(40) <= "00000011010000010101000000100000";
                        f_reg(41) <= "00000001010101000110100000100001";
                        f_reg(42) <= "00101101101100010110111101000101";
                        f_reg(43) <= "00000000110111010111100000000111";
                        f_reg(44) <= "00000010010011110011100000100100";
                        f_reg(45) <= "00000000010100011000000000100101";
                        f_reg(46) <= "00000010110100000010100000100110";
                        f_reg(47) <= "00101110110011100011000111001011";
                        f_reg(48) <= "00101001000000111100000010111011";
                        f_reg(49) <= "00000000101001101110000000100001";
                        f_reg(50) <= "00000011011011001010100000100110";
                        f_reg(51) <= "00000010101111101011100000101011";
                        f_reg(52) <= "00000000000000000000000000000000";
                        f_reg(53) <= "00000000111001001100000000000111";
                        f_reg(54) <= "10101100000010000000010000011100";
                        f_reg(55) <= "00000001011011101001100000100110";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000111101000111000010";
                        f_reg(58) <= "00000000000111000000111001000011";
                        f_reg(59) <= "00100110111010101001000110111000";
                        f_reg(60) <= "10101100000110010000010000100000";
                        f_reg(61) <= "00110100101101001111111000101001";
                        f_reg(62) <= "00100011010011010010111110011100";
                        f_reg(63) <= "00000001001101001110100000100001";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000011000000001001000000101011";
                        f_reg(66) <= "00000011101000010111100000100101";
                        f_reg(67) <= "00000000000000000000000000000000";
                        f_reg(68) <= "00000001010011110001000000100111";
                        f_reg(69) <= "10101100000011010000010000100100";
                        f_reg(70) <= "10101100000100100000010000101000";
                        f_reg(71) <= "10101100000100110000010000101100";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "10101100000000100000010000110000";
                        f_reg(74) <= "00100011111111111111111111111111";
                        f_reg(75) <= "00011111111000001111111110111000";
                        f_reg(76) <= "00010000000000000000000110111101";
                        f_reg(77) <= "00111100000111100000001111100111";
                        f_reg(78) <= "00111100000111110000001111100111";
                        f_reg(79) <= "00000000000111101111010000000010";
                        f_reg(80) <= "00000000000111111111110000000010";
                        f_reg(81) <= "00111100000000011110001011000110";
                        f_reg(82) <= "00111100000011111110001011000110";
                        f_reg(83) <= "00000000000000010001000000100011";
                        f_reg(84) <= "00000000000011111000000000100011";
                        f_reg(85) <= "00110000010000110010110010110100";
                        f_reg(86) <= "00110010000100010010110010110100";
                        f_reg(87) <= "00000000000000100010010111000011";
                        f_reg(88) <= "00000000000100001001010111000011";
                        f_reg(89) <= "00000000100000110010100000100101";
                        f_reg(90) <= "00000010010100011001100000100101";
                        f_reg(91) <= "00000000101001000011000000100111";
                        f_reg(92) <= "00000010011100101010000000100111";
                        f_reg(93) <= "00000000000001000011100000100000";
                        f_reg(94) <= "00000000000100101010100000100000";
                        f_reg(95) <= "00000000110001100100000000100110";
                        f_reg(96) <= "00000010100101001011000000100110";
                        f_reg(97) <= "00000000011001110100100000000110";
                        f_reg(98) <= "00000010001101011011100000000110";
                        f_reg(99) <= "00000000100001010101000000101011";
                        f_reg(100) <= "00000010010100111100000000101011";
                        f_reg(101) <= "00111100000010111011000100000110";
                        f_reg(102) <= "00111100000110011011000100000110";
                        f_reg(103) <= "00000000001000000110000000100111";
                        f_reg(104) <= "00000001111000001101000000100111";
                        f_reg(105) <= "00000000000000000000000000000000";
                        f_reg(106) <= "00000000000000000000000000000000";
                        f_reg(107) <= "00000000100010110110100000100001";
                        f_reg(108) <= "00000010010110011101100000100001";
                        f_reg(109) <= "00000000100000100111000000100100";
                        f_reg(110) <= "00000010010100001110000000100100";
                        f_reg(111) <= "00000001110010010011000000000111";
                        f_reg(112) <= "00000011100101111010000000000111";
                        f_reg(113) <= "00000000000010100000110101000011";
                        f_reg(114) <= "00000000000110000111110101000011";
                        f_reg(115) <= "00000001110010010001000000100110";
                        f_reg(116) <= "00000011100101111000000000100110";
                        f_reg(117) <= "00000001010011010100100000100001";
                        f_reg(118) <= "00000011000110111011100000100001";
                        f_reg(119) <= "00111100000010101111100001001000";
                        f_reg(120) <= "00111100000110001111100001001000";
                        f_reg(121) <= "00110000100011010010101000100001";
                        f_reg(122) <= "00110010010110110010101000100001";
                        f_reg(123) <= "00010101011110010000000100000001";
                        f_reg(124) <= "10101100000010110000010000110100";
                        f_reg(125) <= "00110000010010111110100101000110";
                        f_reg(126) <= "00110010000110011110100101000110";
                        f_reg(127) <= "00000000000001000010010101000011";
                        f_reg(128) <= "00000000000100101001010101000011";
                        f_reg(129) <= "10001100000000100000010000110100";
                        f_reg(130) <= "10001100000100000000010000110100";
                        f_reg(131) <= "00010100010100001111111111111110";
                        f_reg(132) <= "00010101000101100000000011111000";
                        f_reg(133) <= "10101100000010000000010000110100";
                        f_reg(134) <= "00110000010010000000001011101110";
                        f_reg(135) <= "00110010000101100000001011101110";
                        f_reg(136) <= "00010100010100000000000011110100";
                        f_reg(137) <= "10101100000000100000010000111000";
                        f_reg(138) <= "00000000110001110001000000100011";
                        f_reg(139) <= "00000010100101011000000000100011";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000000000000000000000000000";
                        f_reg(142) <= "00000000001000110011000000100010";
                        f_reg(143) <= "00000001111100011010000000100010";
                        f_reg(144) <= "00000001011000100011100000100101";
                        f_reg(145) <= "00000011001100001010100000100101";
                        f_reg(146) <= "00000001110010010000100000100111";
                        f_reg(147) <= "00000011100101110111100000100111";
                        f_reg(148) <= "00010100111101010000000011101000";
                        f_reg(149) <= "10101100000001110000010000111100";
                        f_reg(150) <= "00000000101011100011100000100101";
                        f_reg(151) <= "00000010011111001010100000100101";
                        f_reg(152) <= "10001100000001010000010000111100";
                        f_reg(153) <= "10001100000100110000010000111100";
                        f_reg(154) <= "00010100101100111111111111111110";
                        f_reg(155) <= "00000000101000110111000000000110";
                        f_reg(156) <= "00000010011100011110000000000110";
                        f_reg(157) <= "00110001110000110110101000011011";
                        f_reg(158) <= "00110011100100010110101000011011";
                        f_reg(159) <= "00000001011000100111000000100101";
                        f_reg(160) <= "00000011001100001110000000100101";
                        f_reg(161) <= "00100000110010111011100111011001";
                        f_reg(162) <= "00100010100110011011100111011001";
                        f_reg(163) <= "00000000000010100001010101000011";
                        f_reg(164) <= "00000000000110001000010101000011";
                        f_reg(165) <= "00111100000001101011111011010101";
                        f_reg(166) <= "00111100000101001011111011010101";
                        f_reg(167) <= "10001100000010100000010000111000";
                        f_reg(168) <= "10001100000110000000010000111000";
                        f_reg(169) <= "00010101010110001111111111111110";
                        f_reg(170) <= "00010100101100110000000011010010";
                        f_reg(171) <= "10101100000001010000010000111000";
                        f_reg(172) <= "00000001010001110010100000100101";
                        f_reg(173) <= "00000011000101011001100000100101";
                        f_reg(174) <= "00010100101100110000000011001110";
                        f_reg(175) <= "10101100000001010000010000111100";
                        f_reg(176) <= "00000000001000100010100000100000";
                        f_reg(177) <= "00000001111100001001100000100000";
                        f_reg(178) <= "00000000101011010000100000100001";
                        f_reg(179) <= "00000010011110110111100000100001";
                        f_reg(180) <= "00101100001000100110111101000101";
                        f_reg(181) <= "00101101111100000110111101000101";
                        f_reg(182) <= "00000001011000110010100000000111";
                        f_reg(183) <= "00000011001100011001100000000111";
                        f_reg(184) <= "00000001001001010110100000100100";
                        f_reg(185) <= "00000010111100111101100000100100";
                        f_reg(186) <= "00000000110000100000100000100101";
                        f_reg(187) <= "00000010100100000111100000100101";
                        f_reg(188) <= "00000001000000010001100000100110";
                        f_reg(189) <= "00000010110011111000100000100110";
                        f_reg(190) <= "00101101000010010011000111001011";
                        f_reg(191) <= "00101110110101110011000111001011";
                        f_reg(192) <= "10001100000001010000010000110100";
                        f_reg(193) <= "10001100000100110000010000110100";
                        f_reg(194) <= "00010100101100111111111111111110";
                        f_reg(195) <= "00101000101001101100000010111011";
                        f_reg(196) <= "00101010011101001100000010111011";
                        f_reg(197) <= "00000000011010110001000000100001";
                        f_reg(198) <= "00000010001110011000000000100001";
                        f_reg(199) <= "00000000111011000000100000100110";
                        f_reg(200) <= "00000010101110100111100000100110";
                        f_reg(201) <= "00000000001011100100000000101011";
                        f_reg(202) <= "00000001111111001011000000101011";
                        f_reg(203) <= "00000000000000000000000000000000";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000001101001000101100000000111";
                        f_reg(206) <= "00000011011100101100100000000111";
                        f_reg(207) <= "00010100101100110000000010101101";
                        f_reg(208) <= "10101100000001010000010000011100";
                        f_reg(209) <= "00000001010010010011100000100110";
                        f_reg(210) <= "00000011000101111010100000100110";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000001100110000111000010";
                        f_reg(214) <= "00000000000101001101000111000010";
                        f_reg(215) <= "00000000000000100000111001000011";
                        f_reg(216) <= "00000000000100000111111001000011";
                        f_reg(217) <= "00100101000011101001000110111000";
                        f_reg(218) <= "00100110110111001001000110111000";
                        f_reg(219) <= "10001100000001000000010000111000";
                        f_reg(220) <= "10001100000100100000010000111000";
                        f_reg(221) <= "00010100100100101111111111111110";
                        f_reg(222) <= "00010100100100100000000010011110";
                        f_reg(223) <= "10101100000001000000010000100000";
                        f_reg(224) <= "00110100011011011111111000101001";
                        f_reg(225) <= "00110110001110111111111000101001";
                        f_reg(226) <= "00100001100001010010111110011100";
                        f_reg(227) <= "00100011010100110010111110011100";
                        f_reg(228) <= "10001100000010100000010000111100";
                        f_reg(229) <= "10001100000110000000010000111100";
                        f_reg(230) <= "00010101010110001111111111111110";
                        f_reg(231) <= "00000001010011010100100000100001";
                        f_reg(232) <= "00000011000110111011100000100001";
                        f_reg(233) <= "00000000000000000000000000000000";
                        f_reg(234) <= "00000000000000000000000000000000";
                        f_reg(235) <= "00000001011000000011000000101011";
                        f_reg(236) <= "00000011001000001010000000101011";
                        f_reg(237) <= "00000001001000010001000000100101";
                        f_reg(238) <= "00000010111011111000000000100101";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000001110000100100000000100111";
                        f_reg(242) <= "00000011100100001011000000100111";
                        f_reg(243) <= "00010100101100110000000010001001";
                        f_reg(244) <= "10101100000001010000010000100100";
                        f_reg(245) <= "00010100110101000000000010000111";
                        f_reg(246) <= "10101100000001100000010000101000";
                        f_reg(247) <= "00010100111101010000000010000101";
                        f_reg(248) <= "10101100000001110000010000101100";
                        f_reg(249) <= "00000000000000000000000000000000";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00010101000101100000000010000001";
                        f_reg(252) <= "10101100000010000000010000110000";
                        f_reg(253) <= "00100011110111011111111100000110";
                        f_reg(254) <= "00010011101000000000000000010011";
                        f_reg(255) <= "00100011110111011111111000001100";
                        f_reg(256) <= "00010011101000000000000000010001";
                        f_reg(257) <= "00100011110111011111110100010010";
                        f_reg(258) <= "00010011101000000000000000001111";
                        f_reg(259) <= "00100011110111101111111111111111";
                        f_reg(260) <= "00100011111111111111111111111111";
                        f_reg(261) <= "00010111110111110000000001110111";
                        f_reg(262) <= "00011111111000001111111101001011";
                        f_reg(263) <= "00010000000000000000000100000010";
                        f_reg(264) <= "00000000000000000000000000000000";
                        f_reg(265) <= "00000000000000000000000000000000";
                        f_reg(266) <= "00000000000000000000000000000000";
                        f_reg(267) <= "00000000000000000000000000000000";
                        f_reg(268) <= "00000000000000000000000000000000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "10001100000111010000011110010100";
                        f_reg(274) <= "00011111101000000000000000000011";
                        f_reg(275) <= "00100000000111010000000000111100";
                        f_reg(276) <= "00010000000000000000000000000010";
                        f_reg(277) <= "00100000000111010000000000000000";
                        f_reg(278) <= "00010100001011110000000001100110";
                        f_reg(279) <= "10101111101000010000011100011100";
                        f_reg(280) <= "10001100000111010000011110010100";
                        f_reg(281) <= "00011111101000000000000000000011";
                        f_reg(282) <= "00100000000111010000000000111100";
                        f_reg(283) <= "00010000000000000000000000000010";
                        f_reg(284) <= "00100000000111010000000000000000";
                        f_reg(285) <= "00010100010100000000000001011111";
                        f_reg(286) <= "10101111101000100000011100100000";
                        f_reg(287) <= "10001100000111010000011110010100";
                        f_reg(288) <= "00011111101000000000000000000011";
                        f_reg(289) <= "00100000000111010000000000111100";
                        f_reg(290) <= "00010000000000000000000000000010";
                        f_reg(291) <= "00100000000111010000000000000000";
                        f_reg(292) <= "00010100011100010000000001011000";
                        f_reg(293) <= "10101111101000110000011100100100";
                        f_reg(294) <= "10001100000111010000011110010100";
                        f_reg(295) <= "00011111101000000000000000000011";
                        f_reg(296) <= "00100000000111010000000000111100";
                        f_reg(297) <= "00010000000000000000000000000010";
                        f_reg(298) <= "00100000000111010000000000000000";
                        f_reg(299) <= "00010100100100100000000001010001";
                        f_reg(300) <= "10101111101001000000011100101000";
                        f_reg(301) <= "10001100000111010000011110010100";
                        f_reg(302) <= "00011111101000000000000000000011";
                        f_reg(303) <= "00100000000111010000000000111100";
                        f_reg(304) <= "00010000000000000000000000000010";
                        f_reg(305) <= "00100000000111010000000000000000";
                        f_reg(306) <= "00010100101100110000000001001010";
                        f_reg(307) <= "10101111101001010000011100101100";
                        f_reg(308) <= "10001100000111010000011110010100";
                        f_reg(309) <= "00011111101000000000000000000011";
                        f_reg(310) <= "00100000000111010000000000111100";
                        f_reg(311) <= "00010000000000000000000000000010";
                        f_reg(312) <= "00100000000111010000000000000000";
                        f_reg(313) <= "00010100110101000000000001000011";
                        f_reg(314) <= "10101111101001100000011100110000";
                        f_reg(315) <= "10001100000111010000011110010100";
                        f_reg(316) <= "00011111101000000000000000000011";
                        f_reg(317) <= "00100000000111010000000000111100";
                        f_reg(318) <= "00010000000000000000000000000010";
                        f_reg(319) <= "00100000000111010000000000000000";
                        f_reg(320) <= "00010100111101010000000000111100";
                        f_reg(321) <= "10101111101001110000011100110100";
                        f_reg(322) <= "10001100000111010000011110010100";
                        f_reg(323) <= "00011111101000000000000000000011";
                        f_reg(324) <= "00100000000111010000000000111100";
                        f_reg(325) <= "00010000000000000000000000000010";
                        f_reg(326) <= "00100000000111010000000000000000";
                        f_reg(327) <= "00010101000101100000000000110101";
                        f_reg(328) <= "10101111101010000000011100111000";
                        f_reg(329) <= "10001100000111010000011110010100";
                        f_reg(330) <= "00011111101000000000000000000011";
                        f_reg(331) <= "00100000000111010000000000111100";
                        f_reg(332) <= "00010000000000000000000000000010";
                        f_reg(333) <= "00100000000111010000000000000000";
                        f_reg(334) <= "00010101001101110000000000101110";
                        f_reg(335) <= "10101111101010010000011100111100";
                        f_reg(336) <= "10001100000111010000011110010100";
                        f_reg(337) <= "00011111101000000000000000000011";
                        f_reg(338) <= "00100000000111010000000000111100";
                        f_reg(339) <= "00010000000000000000000000000010";
                        f_reg(340) <= "00100000000111010000000000000000";
                        f_reg(341) <= "00010101010110000000000000100111";
                        f_reg(342) <= "10101111101010100000011101000000";
                        f_reg(343) <= "10001100000111010000011110010100";
                        f_reg(344) <= "00011111101000000000000000000011";
                        f_reg(345) <= "00100000000111010000000000111100";
                        f_reg(346) <= "00010000000000000000000000000010";
                        f_reg(347) <= "00100000000111010000000000000000";
                        f_reg(348) <= "00010101011110010000000000100000";
                        f_reg(349) <= "10101111101010110000011101000100";
                        f_reg(350) <= "10001100000111010000011110010100";
                        f_reg(351) <= "00011111101000000000000000000011";
                        f_reg(352) <= "00100000000111010000000000111100";
                        f_reg(353) <= "00010000000000000000000000000010";
                        f_reg(354) <= "00100000000111010000000000000000";
                        f_reg(355) <= "00010101100110100000000000011001";
                        f_reg(356) <= "10101111101011000000011101001000";
                        f_reg(357) <= "10001100000111010000011110010100";
                        f_reg(358) <= "00011111101000000000000000000011";
                        f_reg(359) <= "00100000000111010000000000111100";
                        f_reg(360) <= "00010000000000000000000000000010";
                        f_reg(361) <= "00100000000111010000000000000000";
                        f_reg(362) <= "00010101101110110000000000010010";
                        f_reg(363) <= "10101111101011010000011101001100";
                        f_reg(364) <= "10001100000111010000011110010100";
                        f_reg(365) <= "00011111101000000000000000000011";
                        f_reg(366) <= "00100000000111010000000000111100";
                        f_reg(367) <= "00010000000000000000000000000010";
                        f_reg(368) <= "00100000000111010000000000000000";
                        f_reg(369) <= "00010101110111000000000000001011";
                        f_reg(370) <= "10101111101011100000011101010000";
                        f_reg(371) <= "10001100000111010000011110010100";
                        f_reg(372) <= "00011111101000000000000000000011";
                        f_reg(373) <= "00100000000111010000000000111100";
                        f_reg(374) <= "00010000000000000000000000000010";
                        f_reg(375) <= "00100000000111010000000000000000";
                        f_reg(376) <= "00010111110111110000000000000100";
                        f_reg(377) <= "10101111101111100000011101010100";
                        f_reg(378) <= "10101100000111010000011110010100";
                        f_reg(379) <= "00010000000000001111111110001000";
                        f_reg(380) <= "10001100000111010000011110010100";
                        f_reg(381) <= "10001111101000010000011100011100";
                        f_reg(382) <= "10001100000111010000011110010100";
                        f_reg(383) <= "10001111101011110000011100011100";
                        f_reg(384) <= "00010100001011111111111111111100";
                        f_reg(385) <= "10001100000111010000011110010100";
                        f_reg(386) <= "10001111101000100000011100100000";
                        f_reg(387) <= "10001100000111010000011110010100";
                        f_reg(388) <= "10001111101100000000011100100000";
                        f_reg(389) <= "00010100010100001111111111111100";
                        f_reg(390) <= "10001100000111010000011110010100";
                        f_reg(391) <= "10001111101000110000011100100100";
                        f_reg(392) <= "10001100000111010000011110010100";
                        f_reg(393) <= "10001111101100010000011100100100";
                        f_reg(394) <= "00010100011100011111111111111100";
                        f_reg(395) <= "10001100000111010000011110010100";
                        f_reg(396) <= "10001111101001000000011100101000";
                        f_reg(397) <= "10001100000111010000011110010100";
                        f_reg(398) <= "10001111101100100000011100101000";
                        f_reg(399) <= "00010100100100101111111111111100";
                        f_reg(400) <= "10001100000111010000011110010100";
                        f_reg(401) <= "10001111101001010000011100101100";
                        f_reg(402) <= "10001100000111010000011110010100";
                        f_reg(403) <= "10001111101100110000011100101100";
                        f_reg(404) <= "00010100101100111111111111111100";
                        f_reg(405) <= "10001100000111010000011110010100";
                        f_reg(406) <= "10001111101001100000011100110000";
                        f_reg(407) <= "10001100000111010000011110010100";
                        f_reg(408) <= "10001111101101000000011100110000";
                        f_reg(409) <= "00010100110101001111111111111100";
                        f_reg(410) <= "10001100000111010000011110010100";
                        f_reg(411) <= "10001111101001110000011100110100";
                        f_reg(412) <= "10001100000111010000011110010100";
                        f_reg(413) <= "10001111101101010000011100110100";
                        f_reg(414) <= "00010100111101011111111111111100";
                        f_reg(415) <= "10001100000111010000011110010100";
                        f_reg(416) <= "10001111101010000000011100111000";
                        f_reg(417) <= "10001100000111010000011110010100";
                        f_reg(418) <= "10001111101101100000011100111000";
                        f_reg(419) <= "00010101000101101111111111111100";
                        f_reg(420) <= "10001100000111010000011110010100";
                        f_reg(421) <= "10001111101010010000011100111100";
                        f_reg(422) <= "10001100000111010000011110010100";
                        f_reg(423) <= "10001111101101110000011100111100";
                        f_reg(424) <= "00010101001101111111111111111100";
                        f_reg(425) <= "10001100000111010000011110010100";
                        f_reg(426) <= "10001111101010100000011101000000";
                        f_reg(427) <= "10001100000111010000011110010100";
                        f_reg(428) <= "10001111101110000000011101000000";
                        f_reg(429) <= "00010101010110001111111111111100";
                        f_reg(430) <= "10001100000111010000011110010100";
                        f_reg(431) <= "10001111101010110000011101000100";
                        f_reg(432) <= "10001100000111010000011110010100";
                        f_reg(433) <= "10001111101110010000011101000100";
                        f_reg(434) <= "00010101011110011111111111111100";
                        f_reg(435) <= "10001100000111010000011110010100";
                        f_reg(436) <= "10001111101011000000011101001000";
                        f_reg(437) <= "10001100000111010000011110010100";
                        f_reg(438) <= "10001111101110100000011101001000";
                        f_reg(439) <= "00010101100110101111111111111100";
                        f_reg(440) <= "10001100000111010000011110010100";
                        f_reg(441) <= "10001111101011010000011101001100";
                        f_reg(442) <= "10001100000111010000011110010100";
                        f_reg(443) <= "10001111101110110000011101001100";
                        f_reg(444) <= "00010101101110111111111111111100";
                        f_reg(445) <= "10001100000111010000011110010100";
                        f_reg(446) <= "10001111101011100000011101010000";
                        f_reg(447) <= "10001100000111010000011110010100";
                        f_reg(448) <= "10001111101111000000011101010000";
                        f_reg(449) <= "00010101110111001111111111111100";
                        f_reg(450) <= "10001100000111010000011110010100";
                        f_reg(451) <= "10001111101111100000011101010100";
                        f_reg(452) <= "10001100000111010000011110010100";
                        f_reg(453) <= "10001111101111110000011101010100";
                        f_reg(454) <= "00010111110111111111111111111100";
                        f_reg(455) <= "00010000000000001111111100111100";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000001111100111";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 -7482
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SUBU R2 R0 R1
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- ANDI R3 R2 11444
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SRA R4 R2 23
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- OR R5 R4 R3
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- NOR R6 R5 R4
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- ADD R7 R0 R4
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- XOR R8 R6 R6
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- SRLV R9 R7 R3
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- SLTU R10 R4 R5
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- LUI R11 -20218
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- NOR R12 R1 R0
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- NOP
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- ADDU R13 R4 R11
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- AND R14 R4 R2
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- SRAV R15 R9 R14
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SRA R16 R10 21
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- XOR R17 R14 R9
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- ADDU R18 R10 R13
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- LUI R19 -1976
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- ANDI R20 R4 10785
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- ANDI R21 R17 -5818
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- SRA R4 R4 21
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- ANDI R22 R11 750
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- SUBU R23 R15 R7
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- NOP
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- SUB R24 R16 R3
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- OR R25 R21 R23
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- NOR R26 R14 R18
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- OR R27 R5 R14
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- SRLV R28 R3 R25
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- ANDI R29 R28 27163
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- OR R30 R21 R23
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- ADDI R6 R24 -17959
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- SRA R1 R19 21
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- LUI R2 -16683
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- OR R9 R11 R27
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- ADD R10 R26 R1
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- ADDU R13 R10 R20
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- SLTIU R17 R13 28485
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SRAV R15 R29 R6
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- AND R7 R18 R15
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- OR R16 R2 R17
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- XOR R5 R22 R16
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- SLTIU R14 R22 12747
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- SLTI R3 R8 -16197
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- ADDU R28 R5 R6
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- XOR R21 R27 R12
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SLTU R23 R21 R30
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- NOP
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- SRAV R24 R4 R7
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SW R8 R0 1052
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- XOR R19 R11 R14
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- NOP
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SRL R26 R3 7
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- SRA R1 R28 25
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- ADDIU R10 R23 -28232
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SW R25 R0 1056
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- ORI R20 R5 -471
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- ADDI R13 R26 12188
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- ADDU R29 R9 R20
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- NOP
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- SLTU R18 R24 R0
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- OR R15 R29 R1
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- NOP
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- NOR R2 R10 R15
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- SW R13 R0 1060
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SW R18 R0 1064
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- SW R19 R0 1068
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- NOP
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SW R2 R0 1072
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- ADDI R31 R31 -1
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- BGTZ R31 -72
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- BEQ R0 R0 445
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- LUI R30 999
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- LUI R31 999
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- SRL R30 R30 16
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- SRL R31 R31 16
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- LUI R1 -7482
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- LUI R15 -7482
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SUBU R2 R0 R1
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- SUBU R16 R0 R15
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- ANDI R3 R2 11444
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- ANDI R17 R16 11444
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SRA R4 R2 23
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- SRA R18 R16 23
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- OR R5 R4 R3
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- OR R19 R18 R17
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- NOR R6 R5 R4
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- NOR R20 R19 R18
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- ADD R7 R0 R4
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- ADD R21 R0 R18
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- XOR R8 R6 R6
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- XOR R22 R20 R20
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SRLV R9 R7 R3
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SRLV R23 R21 R17
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- SLTU R10 R4 R5
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- SLTU R24 R18 R19
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- LUI R11 -20218
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- LUI R25 -20218
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- NOR R12 R1 R0
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- NOR R26 R15 R0
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- NOP
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- NOP
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- ADDU R13 R4 R11
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- ADDU R27 R18 R25
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- AND R14 R4 R2
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- AND R28 R18 R16
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- SRAV R6 R9 R14
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- SRAV R20 R23 R28
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- SRA R1 R10 21
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- SRA R15 R24 21
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- XOR R2 R14 R9
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- XOR R16 R28 R23
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- ADDU R9 R10 R13
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- ADDU R23 R24 R27
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- LUI R10 -1976
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- LUI R24 -1976
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- ANDI R13 R4 10785
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- ANDI R27 R18 10785
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- BNE R11 R25 257
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SW R11 R0 1076
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- ANDI R11 R2 -5818
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- ANDI R25 R16 -5818
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- SRA R4 R4 21
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SRA R18 R18 21
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- LW R2 R0 1076
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- LW R16 R0 1076
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- BNE R2 R16 -2
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- BNE R8 R22 248
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- SW R8 R0 1076
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- ANDI R8 R2 750
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- ANDI R22 R16 750
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- BNE R2 R16 244
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- SW R2 R0 1080
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SUBU R2 R6 R7
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- SUBU R16 R20 R21
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- NOP
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- NOP
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- SUB R6 R1 R3
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- SUB R20 R15 R17
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- OR R7 R11 R2
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- OR R21 R25 R16
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- NOR R1 R14 R9
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- NOR R15 R28 R23
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- BNE R7 R21 232
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- SW R7 R0 1084
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- OR R7 R5 R14
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- OR R21 R19 R28
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- LW R5 R0 1084
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- LW R19 R0 1084
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- BNE R5 R19 -2
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- SRLV R14 R3 R5
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- SRLV R28 R17 R19
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- ANDI R3 R14 27163
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- ANDI R17 R28 27163
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- OR R14 R11 R2
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- OR R28 R25 R16
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- ADDI R11 R6 -17959
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- ADDI R25 R20 -17959
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- SRA R2 R10 21
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- SRA R16 R24 21
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- LUI R6 -16683
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- LUI R20 -16683
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- LW R10 R0 1080
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- LW R24 R0 1080
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- BNE R10 R24 -2
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- BNE R5 R19 210
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- SW R5 R0 1080
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- OR R5 R10 R7
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- OR R19 R24 R21
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- BNE R5 R19 206
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- SW R5 R0 1084
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- ADD R5 R1 R2
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- ADD R19 R15 R16
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- ADDU R1 R5 R13
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- ADDU R15 R19 R27
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- SLTIU R2 R1 28485
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- SLTIU R16 R15 28485
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SRAV R5 R3 R11
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- SRAV R19 R17 R25
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- AND R13 R9 R5
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- AND R27 R23 R19
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- OR R1 R6 R2
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- OR R15 R20 R16
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- XOR R3 R8 R1
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- XOR R17 R22 R15
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- SLTIU R9 R8 12747
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- SLTIU R23 R22 12747
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- LW R5 R0 1076
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- LW R19 R0 1076
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- BNE R5 R19 -2
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- SLTI R6 R5 -16197
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- SLTI R20 R19 -16197
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- ADDU R2 R3 R11
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- ADDU R16 R17 R25
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- XOR R1 R7 R12
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- XOR R15 R21 R26
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- SLTU R8 R1 R14
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- SLTU R22 R15 R28
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- NOP
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- NOP
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- SRAV R11 R4 R13
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- SRAV R25 R18 R27
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- BNE R5 R19 173
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- SW R5 R0 1052
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- XOR R7 R10 R9
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- XOR R21 R24 R23
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- NOP
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- NOP
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- SRL R12 R6 7
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- SRL R26 R20 7
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- SRA R1 R2 25
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- SRA R15 R16 25
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- ADDIU R14 R8 -28232
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- ADDIU R28 R22 -28232
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- LW R4 R0 1080
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- LW R18 R0 1080
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- BNE R4 R18 -2
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- BNE R4 R18 158
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- SW R4 R0 1056
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- ORI R13 R3 -471
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- ORI R27 R17 -471
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- ADDI R5 R12 12188
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- ADDI R19 R26 12188
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- LW R10 R0 1084
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- LW R24 R0 1084
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- BNE R10 R24 -2
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- ADDU R9 R10 R13
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- ADDU R23 R24 R27
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- NOP
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- NOP
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- SLTU R6 R11 R0
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- SLTU R20 R25 R0
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- OR R2 R9 R1
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- OR R16 R23 R15
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- NOP
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- NOP
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- NOR R8 R14 R2
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- NOR R22 R28 R16
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- BNE R5 R19 137
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- SW R5 R0 1060
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- BNE R6 R20 135
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- SW R6 R0 1064
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- BNE R7 R21 133
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- SW R7 R0 1068
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- NOP
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- NOP
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- BNE R8 R22 129
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- SW R8 R0 1072
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- ADDI R29 R30 -250
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- BEQ R29 R0 19
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- ADDI R29 R30 -500
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- BEQ R29 R0 17
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- ADDI R29 R30 -750
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- BEQ R29 R0 15
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- ADDI R30 R30 -1
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- ADDI R31 R31 -1
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- BNE R30 R31 119
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- BGTZ R31 -181
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- BEQ R0 R0 258
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- NOP
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- NOP
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- NOP
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- NOP
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- NOP
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- NOP
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- NOP
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- NOP
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- NOP
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- LW R29 R0 1940
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- BGTZ R29 3
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- ADDI R29 R0 60
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- BEQ R0 R0 2
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- ADDI R29 R0 0
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- BNE R1 R15 102
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- SW R1 R29 1820
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- LW R29 R0 1940
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- BGTZ R29 3
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- ADDI R29 R0 60
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- BEQ R0 R0 2
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- ADDI R29 R0 0
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- BNE R2 R16 95
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- SW R2 R29 1824
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- LW R29 R0 1940
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- BGTZ R29 3
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- ADDI R29 R0 60
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- BEQ R0 R0 2
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- ADDI R29 R0 0
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- BNE R3 R17 88
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- SW R3 R29 1828
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- LW R29 R0 1940
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- BGTZ R29 3
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- ADDI R29 R0 60
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- BEQ R0 R0 2
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- ADDI R29 R0 0
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- BNE R4 R18 81
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- SW R4 R29 1832
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- LW R29 R0 1940
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- BGTZ R29 3
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- ADDI R29 R0 60
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- BEQ R0 R0 2
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- ADDI R29 R0 0
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- BNE R5 R19 74
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- SW R5 R29 1836
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- LW R29 R0 1940
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- BGTZ R29 3
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- ADDI R29 R0 60
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- BEQ R0 R0 2
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- ADDI R29 R0 0
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- BNE R6 R20 67
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- SW R6 R29 1840
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- LW R29 R0 1940
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- BGTZ R29 3
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- ADDI R29 R0 60
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- BEQ R0 R0 2
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- ADDI R29 R0 0
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- BNE R7 R21 60
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- SW R7 R29 1844
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- LW R29 R0 1940
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- BGTZ R29 3
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- ADDI R29 R0 60
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- BEQ R0 R0 2
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- ADDI R29 R0 0
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- BNE R8 R22 53
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- SW R8 R29 1848
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- LW R29 R0 1940
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- BGTZ R29 3
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- ADDI R29 R0 60
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- BEQ R0 R0 2
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- ADDI R29 R0 0
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- BNE R9 R23 46
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- SW R9 R29 1852
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- LW R29 R0 1940
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- BGTZ R29 3
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- ADDI R29 R0 60
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- BEQ R0 R0 2
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- ADDI R29 R0 0
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- BNE R10 R24 39
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- SW R10 R29 1856
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- LW R29 R0 1940
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- BGTZ R29 3
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- ADDI R29 R0 60
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- BEQ R0 R0 2
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- ADDI R29 R0 0
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- BNE R11 R25 32
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- SW R11 R29 1860
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- LW R29 R0 1940
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- BGTZ R29 3
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- ADDI R29 R0 60
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- BEQ R0 R0 2
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- ADDI R29 R0 0
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- BNE R12 R26 25
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- SW R12 R29 1864
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- LW R29 R0 1940
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- BGTZ R29 3
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- ADDI R29 R0 60
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- BEQ R0 R0 2
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- ADDI R29 R0 0
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- BNE R13 R27 18
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- SW R13 R29 1868
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- LW R29 R0 1940
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- BGTZ R29 3
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- ADDI R29 R0 60
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- BEQ R0 R0 2
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- ADDI R29 R0 0
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- BNE R14 R28 11
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- SW R14 R29 1872
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- LW R29 R0 1940
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- BGTZ R29 3
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- ADDI R29 R0 60
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- BEQ R0 R0 2
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- ADDI R29 R0 0
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- BNE R30 R31 4
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- SW R30 R29 1876
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- SW R29 R0 1940
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- BEQ R0 R0 -120
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- LW R29 R0 1940
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- LW R1 R29 1820
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- LW R29 R0 1940
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- LW R15 R29 1820
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- BNE R1 R15 -4
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- LW R29 R0 1940
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- LW R2 R29 1824
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- LW R29 R0 1940
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- LW R16 R29 1824
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- BNE R2 R16 -4
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- LW R29 R0 1940
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- LW R3 R29 1828
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- LW R29 R0 1940
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- LW R17 R29 1828
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- BNE R3 R17 -4
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- LW R29 R0 1940
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- LW R4 R29 1832
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- LW R29 R0 1940
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- LW R18 R29 1832
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- BNE R4 R18 -4
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- LW R29 R0 1940
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- LW R5 R29 1836
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- LW R29 R0 1940
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- LW R19 R29 1836
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- BNE R5 R19 -4
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- LW R29 R0 1940
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- LW R6 R29 1840
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- LW R29 R0 1940
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- LW R20 R29 1840
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- BNE R6 R20 -4
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- LW R29 R0 1940
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- LW R7 R29 1844
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- LW R29 R0 1940
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- LW R21 R29 1844
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- BNE R7 R21 -4
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- LW R29 R0 1940
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- LW R8 R29 1848
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- LW R29 R0 1940
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- LW R22 R29 1848
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- BNE R8 R22 -4
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- LW R29 R0 1940
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- LW R9 R29 1852
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- LW R29 R0 1940
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- LW R23 R29 1852
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- BNE R9 R23 -4
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R29 R0 1940
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R10 R29 1856
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- LW R29 R0 1940
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- LW R24 R29 1856
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- BNE R10 R24 -4
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- LW R29 R0 1940
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- LW R11 R29 1860
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- LW R29 R0 1940
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- LW R25 R29 1860
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- BNE R11 R25 -4
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- LW R29 R0 1940
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- LW R12 R29 1864
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- LW R29 R0 1940
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- LW R26 R29 1864
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- BNE R12 R26 -4
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- LW R29 R0 1940
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- LW R13 R29 1868
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- LW R29 R0 1940
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- LW R27 R29 1868
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- BNE R13 R27 -4
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- LW R29 R0 1940
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- LW R14 R29 1872
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- LW R29 R0 1940
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- LW R28 R29 1872
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- BNE R14 R28 -4
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- LW R29 R0 1940
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- LW R30 R29 1876
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- LW R29 R0 1940
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- LW R31 R29 1876
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- BNE R30 R31 -4
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- BEQ R0 R0 -196
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- NOP
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- NOP
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- NOP
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- NOP
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- NOP
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- NOP
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- NOP
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- NOP
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- NOP
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- NOP
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- NOP
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- NOP
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- NOP
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- NOP
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- NOP
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- NOP
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- NOP
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- NOP
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- NOP
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- NOP
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- NOP
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- NOP
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- NOP
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- NOP
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- NOP
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- NOP
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- NOP
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- NOP
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- NOP
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- NOP
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- NOP
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- NOP
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- NOP
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- NOP
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- NOP
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- NOP
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- NOP
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- NOP
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- NOP
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- NOP
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- NOP
                        f_reg(496) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(497) =>
                        -- NOP
                        f_reg(497) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(498) =>
                        -- NOP
                        f_reg(498) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(499) =>
                        -- NOP
                        f_reg(499) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(500) =>
                        -- NOP
                        f_reg(500) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(501) =>
                        -- NOP
                        f_reg(501) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(502) =>
                        -- NOP
                        f_reg(502) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(503) =>
                        -- NOP
                        f_reg(503) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(504) =>
                        -- NOP
                        f_reg(504) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(505) =>
                        -- NOP
                        f_reg(505) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(506) =>
                        -- NOP
                        f_reg(506) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(507) =>
                        -- NOP
                        f_reg(507) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(508) =>
                        -- NOP
                        f_reg(508) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(509) =>
                        -- NOP
                        f_reg(509) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(510) =>
                        -- NOP
                        f_reg(510) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(511) =>
                        -- NOP
                        f_reg(511) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(512) =>
                        -- NOP
                        f_reg(512) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(513) =>
                        -- NOP
                        f_reg(513) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(514) =>
                        -- NOP
                        f_reg(514) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(515) =>
                        -- NOP
                        f_reg(515) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(516) =>
                        -- NOP
                        f_reg(516) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(517) =>
                        -- NOP
                        f_reg(517) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(518) =>
                        -- NOP
                        f_reg(518) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(519) =>
                        -- NOP
                        f_reg(519) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(520) =>
                        -- NOP
                        f_reg(520) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(521) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011110001011000110";
                        f_reg(4) <= "00000000000000010001000000100011";
                        f_reg(5) <= "00110000010000110010110010110100";
                        f_reg(6) <= "00000000000000100010010111000011";
                        f_reg(7) <= "00000000100000110010100000100101";
                        f_reg(8) <= "00000000101001000011000000100111";
                        f_reg(9) <= "00000000000001000011100000100000";
                        f_reg(10) <= "00000000110001100100000000100110";
                        f_reg(11) <= "00000000011001110100100000000110";
                        f_reg(12) <= "00000000100001010101000000101011";
                        f_reg(13) <= "00111100000010111011000100000110";
                        f_reg(14) <= "00000000001000000110000000100111";
                        f_reg(15) <= "00000000000000000000000000000000";
                        f_reg(16) <= "00000000100010110110100000100001";
                        f_reg(17) <= "00000000100000100111000000100100";
                        f_reg(18) <= "00000001110010010111100000000111";
                        f_reg(19) <= "00000000000010101000010101000011";
                        f_reg(20) <= "00000001110010011000100000100110";
                        f_reg(21) <= "00000001010011011001000000100001";
                        f_reg(22) <= "00111100000100111111100001001000";
                        f_reg(23) <= "00110000100101000010101000100001";
                        f_reg(24) <= "00110010001101011110100101000110";
                        f_reg(25) <= "00000000000001000010010101000011";
                        f_reg(26) <= "00110001011101100000001011101110";
                        f_reg(27) <= "00000001111001111011100000100011";
                        f_reg(28) <= "00000000000000000000000000000000";
                        f_reg(29) <= "00000010000000111100000000100010";
                        f_reg(30) <= "00000010101101111100100000100101";
                        f_reg(31) <= "00000001110100101101000000100111";
                        f_reg(32) <= "00000000101011101101100000100101";
                        f_reg(33) <= "00000011001000111110000000000110";
                        f_reg(34) <= "00110011100111010110101000011011";
                        f_reg(35) <= "00000010101101111111000000100101";
                        f_reg(36) <= "00100011000001101011100111011001";
                        f_reg(37) <= "00000000000100110000110101000011";
                        f_reg(38) <= "00111100000000101011111011010101";
                        f_reg(39) <= "00000001011110110100100000100101";
                        f_reg(40) <= "00000011010000010101000000100000";
                        f_reg(41) <= "00000001010101000110100000100001";
                        f_reg(42) <= "00101101101100010110111101000101";
                        f_reg(43) <= "00000000110111010111100000000111";
                        f_reg(44) <= "00000010010011110011100000100100";
                        f_reg(45) <= "00000000010100011000000000100101";
                        f_reg(46) <= "00000010110100000010100000100110";
                        f_reg(47) <= "00101110110011100011000111001011";
                        f_reg(48) <= "00101001000000111100000010111011";
                        f_reg(49) <= "00000000101001101110000000100001";
                        f_reg(50) <= "00000011011011001010100000100110";
                        f_reg(51) <= "00000010101111101011100000101011";
                        f_reg(52) <= "00000000000000000000000000000000";
                        f_reg(53) <= "00000000111001001100000000000111";
                        f_reg(54) <= "10101100000010000000010000011100";
                        f_reg(55) <= "00000001011011101001100000100110";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000111101000111000010";
                        f_reg(58) <= "00000000000111000000111001000011";
                        f_reg(59) <= "00100110111010101001000110111000";
                        f_reg(60) <= "10101100000110010000010000100000";
                        f_reg(61) <= "00110100101101001111111000101001";
                        f_reg(62) <= "00100011010011010010111110011100";
                        f_reg(63) <= "00000001001101001110100000100001";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000011000000001001000000101011";
                        f_reg(66) <= "00000011101000010111100000100101";
                        f_reg(67) <= "00000000000000000000000000000000";
                        f_reg(68) <= "00000001010011110001000000100111";
                        f_reg(69) <= "10101100000011010000010000100100";
                        f_reg(70) <= "10101100000100100000010000101000";
                        f_reg(71) <= "10101100000100110000010000101100";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "10101100000000100000010000110000";
                        f_reg(74) <= "00100011111111111111111111111111";
                        f_reg(75) <= "00011111111000001111111110111000";
                        f_reg(76) <= "00010000000000000000000110111101";
                        f_reg(77) <= "00111100000111100000001111100111";
                        f_reg(78) <= "00111100000111110000001111100111";
                        f_reg(79) <= "00000000000111101111010000000010";
                        f_reg(80) <= "00000000000111111111110000000010";
                        f_reg(81) <= "00111100000000011110001011000110";
                        f_reg(82) <= "00111100000011111110001011000110";
                        f_reg(83) <= "00000000000000010001000000100011";
                        f_reg(84) <= "00000000000011111000000000100011";
                        f_reg(85) <= "00110000010000110010110010110100";
                        f_reg(86) <= "00110010000100010010110010110100";
                        f_reg(87) <= "00000000000000100010010111000011";
                        f_reg(88) <= "00000000000100001001010111000011";
                        f_reg(89) <= "00000000100000110010100000100101";
                        f_reg(90) <= "00000010010100011001100000100101";
                        f_reg(91) <= "00000000101001000011000000100111";
                        f_reg(92) <= "00000010011100101010000000100111";
                        f_reg(93) <= "00000000000001000011100000100000";
                        f_reg(94) <= "00000000000100101010100000100000";
                        f_reg(95) <= "00000000110001100100000000100110";
                        f_reg(96) <= "00000010100101001011000000100110";
                        f_reg(97) <= "00000000011001110100100000000110";
                        f_reg(98) <= "00000010001101011011100000000110";
                        f_reg(99) <= "00000000100001010101000000101011";
                        f_reg(100) <= "00000010010100111100000000101011";
                        f_reg(101) <= "00111100000010111011000100000110";
                        f_reg(102) <= "00111100000110011011000100000110";
                        f_reg(103) <= "00000000001000000110000000100111";
                        f_reg(104) <= "00000001111000001101000000100111";
                        f_reg(105) <= "00000000000000000000000000000000";
                        f_reg(106) <= "00000000000000000000000000000000";
                        f_reg(107) <= "00000000100010110110100000100001";
                        f_reg(108) <= "00000010010110011101100000100001";
                        f_reg(109) <= "00000000100000100111000000100100";
                        f_reg(110) <= "00000010010100001110000000100100";
                        f_reg(111) <= "00000001110010010011000000000111";
                        f_reg(112) <= "00000011100101111010000000000111";
                        f_reg(113) <= "00000000000010100000110101000011";
                        f_reg(114) <= "00000000000110000111110101000011";
                        f_reg(115) <= "00000001110010010001000000100110";
                        f_reg(116) <= "00000011100101111000000000100110";
                        f_reg(117) <= "00000001010011010100100000100001";
                        f_reg(118) <= "00000011000110111011100000100001";
                        f_reg(119) <= "00111100000010101111100001001000";
                        f_reg(120) <= "00111100000110001111100001001000";
                        f_reg(121) <= "00110000100011010010101000100001";
                        f_reg(122) <= "00110010010110110010101000100001";
                        f_reg(123) <= "00010101011110010000000100000001";
                        f_reg(124) <= "10101100000010110000010000110100";
                        f_reg(125) <= "00110000010010111110100101000110";
                        f_reg(126) <= "00110010000110011110100101000110";
                        f_reg(127) <= "00000000000001000010010101000011";
                        f_reg(128) <= "00000000000100101001010101000011";
                        f_reg(129) <= "10001100000000100000010000110100";
                        f_reg(130) <= "10001100000100000000010000110100";
                        f_reg(131) <= "00010100010100001111111111111110";
                        f_reg(132) <= "00010101000101100000000011111000";
                        f_reg(133) <= "10101100000010000000010000110100";
                        f_reg(134) <= "00110000010010000000001011101110";
                        f_reg(135) <= "00110010000101100000001011101110";
                        f_reg(136) <= "00010100010100000000000011110100";
                        f_reg(137) <= "10101100000000100000010000111000";
                        f_reg(138) <= "00000000110001110001000000100011";
                        f_reg(139) <= "00000010100101011000000000100011";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000000000000000000000000000";
                        f_reg(142) <= "00000000001000110011000000100010";
                        f_reg(143) <= "00000001111100011010000000100010";
                        f_reg(144) <= "00000001011000100011100000100101";
                        f_reg(145) <= "00000011001100001010100000100101";
                        f_reg(146) <= "00000001110010010000100000100111";
                        f_reg(147) <= "00000011100101110111100000100111";
                        f_reg(148) <= "00010100111101010000000011101000";
                        f_reg(149) <= "10101100000001110000010000111100";
                        f_reg(150) <= "00000000101011100011100000100101";
                        f_reg(151) <= "00000010011111001010100000100101";
                        f_reg(152) <= "10001100000001010000010000111100";
                        f_reg(153) <= "10001100000100110000010000111100";
                        f_reg(154) <= "00010100101100111111111111111110";
                        f_reg(155) <= "00000000101000110111000000000110";
                        f_reg(156) <= "00000010011100011110000000000110";
                        f_reg(157) <= "00110001110000110110101000011011";
                        f_reg(158) <= "00110011100100010110101000011011";
                        f_reg(159) <= "00000001011000100111000000100101";
                        f_reg(160) <= "00000011001100001110000000100101";
                        f_reg(161) <= "00100000110010111011100111011001";
                        f_reg(162) <= "00100010100110011011100111011001";
                        f_reg(163) <= "00000000000010100001010101000011";
                        f_reg(164) <= "00000000000110001000010101000011";
                        f_reg(165) <= "00111100000001101011111011010101";
                        f_reg(166) <= "00111100000101001011111011010101";
                        f_reg(167) <= "10001100000010100000010000111000";
                        f_reg(168) <= "10001100000110000000010000111000";
                        f_reg(169) <= "00010101010110001111111111111110";
                        f_reg(170) <= "00010100101100110000000011010010";
                        f_reg(171) <= "10101100000001010000010000111000";
                        f_reg(172) <= "00000001010001110010100000100101";
                        f_reg(173) <= "00000011000101011001100000100101";
                        f_reg(174) <= "00010100101100110000000011001110";
                        f_reg(175) <= "10101100000001010000010000111100";
                        f_reg(176) <= "00000000001000100010100000100000";
                        f_reg(177) <= "00000001111100001001100000100000";
                        f_reg(178) <= "00000000101011010000100000100001";
                        f_reg(179) <= "00000010011110110111100000100001";
                        f_reg(180) <= "00101100001000100110111101000101";
                        f_reg(181) <= "00101101111100000110111101000101";
                        f_reg(182) <= "00000001011000110010100000000111";
                        f_reg(183) <= "00000011001100011001100000000111";
                        f_reg(184) <= "00000001001001010110100000100100";
                        f_reg(185) <= "00000010111100111101100000100100";
                        f_reg(186) <= "00000000110000100000100000100101";
                        f_reg(187) <= "00000010100100000111100000100101";
                        f_reg(188) <= "00000001000000010001100000100110";
                        f_reg(189) <= "00000010110011111000100000100110";
                        f_reg(190) <= "00101101000010010011000111001011";
                        f_reg(191) <= "00101110110101110011000111001011";
                        f_reg(192) <= "10001100000001010000010000110100";
                        f_reg(193) <= "10001100000100110000010000110100";
                        f_reg(194) <= "00010100101100111111111111111110";
                        f_reg(195) <= "00101000101001101100000010111011";
                        f_reg(196) <= "00101010011101001100000010111011";
                        f_reg(197) <= "00000000011010110001000000100001";
                        f_reg(198) <= "00000010001110011000000000100001";
                        f_reg(199) <= "00000000111011000000100000100110";
                        f_reg(200) <= "00000010101110100111100000100110";
                        f_reg(201) <= "00000000001011100100000000101011";
                        f_reg(202) <= "00000001111111001011000000101011";
                        f_reg(203) <= "00000000000000000000000000000000";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000001101001000101100000000111";
                        f_reg(206) <= "00000011011100101100100000000111";
                        f_reg(207) <= "00010100101100110000000010101101";
                        f_reg(208) <= "10101100000001010000010000011100";
                        f_reg(209) <= "00000001010010010011100000100110";
                        f_reg(210) <= "00000011000101111010100000100110";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000001100110000111000010";
                        f_reg(214) <= "00000000000101001101000111000010";
                        f_reg(215) <= "00000000000000100000111001000011";
                        f_reg(216) <= "00000000000100000111111001000011";
                        f_reg(217) <= "00100101000011101001000110111000";
                        f_reg(218) <= "00100110110111001001000110111000";
                        f_reg(219) <= "10001100000001000000010000111000";
                        f_reg(220) <= "10001100000100100000010000111000";
                        f_reg(221) <= "00010100100100101111111111111110";
                        f_reg(222) <= "00010100100100100000000010011110";
                        f_reg(223) <= "10101100000001000000010000100000";
                        f_reg(224) <= "00110100011011011111111000101001";
                        f_reg(225) <= "00110110001110111111111000101001";
                        f_reg(226) <= "00100001100001010010111110011100";
                        f_reg(227) <= "00100011010100110010111110011100";
                        f_reg(228) <= "10001100000010100000010000111100";
                        f_reg(229) <= "10001100000110000000010000111100";
                        f_reg(230) <= "00010101010110001111111111111110";
                        f_reg(231) <= "00000001010011010100100000100001";
                        f_reg(232) <= "00000011000110111011100000100001";
                        f_reg(233) <= "00000000000000000000000000000000";
                        f_reg(234) <= "00000000000000000000000000000000";
                        f_reg(235) <= "00000001011000000011000000101011";
                        f_reg(236) <= "00000011001000001010000000101011";
                        f_reg(237) <= "00000001001000010001000000100101";
                        f_reg(238) <= "00000010111011111000000000100101";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000001110000100100000000100111";
                        f_reg(242) <= "00000011100100001011000000100111";
                        f_reg(243) <= "00010100101100110000000010001001";
                        f_reg(244) <= "10101100000001010000010000100100";
                        f_reg(245) <= "00010100110101000000000010000111";
                        f_reg(246) <= "10101100000001100000010000101000";
                        f_reg(247) <= "00010100111101010000000010000101";
                        f_reg(248) <= "10101100000001110000010000101100";
                        f_reg(249) <= "00000000000000000000000000000000";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00010101000101100000000010000001";
                        f_reg(252) <= "10101100000010000000010000110000";
                        f_reg(253) <= "00100011110111011111111100000110";
                        f_reg(254) <= "00010011101000000000000000010011";
                        f_reg(255) <= "00100011110111011111111000001100";
                        f_reg(256) <= "00010011101000000000000000010001";
                        f_reg(257) <= "00100011110111011111110100010010";
                        f_reg(258) <= "00010011101000000000000000001111";
                        f_reg(259) <= "00100011110111101111111111111111";
                        f_reg(260) <= "00100011111111111111111111111111";
                        f_reg(261) <= "00010111110111110000000001110111";
                        f_reg(262) <= "00011111111000001111111101001011";
                        f_reg(263) <= "00010000000000000000000100000010";
                        f_reg(264) <= "00000000000000000000000000000000";
                        f_reg(265) <= "00000000000000000000000000000000";
                        f_reg(266) <= "00000000000000000000000000000000";
                        f_reg(267) <= "00000000000000000000000000000000";
                        f_reg(268) <= "00000000000000000000000000000000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "10001100000111010000011110010100";
                        f_reg(274) <= "00011111101000000000000000000011";
                        f_reg(275) <= "00100000000111010000000000111100";
                        f_reg(276) <= "00010000000000000000000000000010";
                        f_reg(277) <= "00100000000111010000000000000000";
                        f_reg(278) <= "00010100001011110000000001100110";
                        f_reg(279) <= "10101111101000010000011100011100";
                        f_reg(280) <= "10001100000111010000011110010100";
                        f_reg(281) <= "00011111101000000000000000000011";
                        f_reg(282) <= "00100000000111010000000000111100";
                        f_reg(283) <= "00010000000000000000000000000010";
                        f_reg(284) <= "00100000000111010000000000000000";
                        f_reg(285) <= "00010100010100000000000001011111";
                        f_reg(286) <= "10101111101000100000011100100000";
                        f_reg(287) <= "10001100000111010000011110010100";
                        f_reg(288) <= "00011111101000000000000000000011";
                        f_reg(289) <= "00100000000111010000000000111100";
                        f_reg(290) <= "00010000000000000000000000000010";
                        f_reg(291) <= "00100000000111010000000000000000";
                        f_reg(292) <= "00010100011100010000000001011000";
                        f_reg(293) <= "10101111101000110000011100100100";
                        f_reg(294) <= "10001100000111010000011110010100";
                        f_reg(295) <= "00011111101000000000000000000011";
                        f_reg(296) <= "00100000000111010000000000111100";
                        f_reg(297) <= "00010000000000000000000000000010";
                        f_reg(298) <= "00100000000111010000000000000000";
                        f_reg(299) <= "00010100100100100000000001010001";
                        f_reg(300) <= "10101111101001000000011100101000";
                        f_reg(301) <= "10001100000111010000011110010100";
                        f_reg(302) <= "00011111101000000000000000000011";
                        f_reg(303) <= "00100000000111010000000000111100";
                        f_reg(304) <= "00010000000000000000000000000010";
                        f_reg(305) <= "00100000000111010000000000000000";
                        f_reg(306) <= "00010100101100110000000001001010";
                        f_reg(307) <= "10101111101001010000011100101100";
                        f_reg(308) <= "10001100000111010000011110010100";
                        f_reg(309) <= "00011111101000000000000000000011";
                        f_reg(310) <= "00100000000111010000000000111100";
                        f_reg(311) <= "00010000000000000000000000000010";
                        f_reg(312) <= "00100000000111010000000000000000";
                        f_reg(313) <= "00010100110101000000000001000011";
                        f_reg(314) <= "10101111101001100000011100110000";
                        f_reg(315) <= "10001100000111010000011110010100";
                        f_reg(316) <= "00011111101000000000000000000011";
                        f_reg(317) <= "00100000000111010000000000111100";
                        f_reg(318) <= "00010000000000000000000000000010";
                        f_reg(319) <= "00100000000111010000000000000000";
                        f_reg(320) <= "00010100111101010000000000111100";
                        f_reg(321) <= "10101111101001110000011100110100";
                        f_reg(322) <= "10001100000111010000011110010100";
                        f_reg(323) <= "00011111101000000000000000000011";
                        f_reg(324) <= "00100000000111010000000000111100";
                        f_reg(325) <= "00010000000000000000000000000010";
                        f_reg(326) <= "00100000000111010000000000000000";
                        f_reg(327) <= "00010101000101100000000000110101";
                        f_reg(328) <= "10101111101010000000011100111000";
                        f_reg(329) <= "10001100000111010000011110010100";
                        f_reg(330) <= "00011111101000000000000000000011";
                        f_reg(331) <= "00100000000111010000000000111100";
                        f_reg(332) <= "00010000000000000000000000000010";
                        f_reg(333) <= "00100000000111010000000000000000";
                        f_reg(334) <= "00010101001101110000000000101110";
                        f_reg(335) <= "10101111101010010000011100111100";
                        f_reg(336) <= "10001100000111010000011110010100";
                        f_reg(337) <= "00011111101000000000000000000011";
                        f_reg(338) <= "00100000000111010000000000111100";
                        f_reg(339) <= "00010000000000000000000000000010";
                        f_reg(340) <= "00100000000111010000000000000000";
                        f_reg(341) <= "00010101010110000000000000100111";
                        f_reg(342) <= "10101111101010100000011101000000";
                        f_reg(343) <= "10001100000111010000011110010100";
                        f_reg(344) <= "00011111101000000000000000000011";
                        f_reg(345) <= "00100000000111010000000000111100";
                        f_reg(346) <= "00010000000000000000000000000010";
                        f_reg(347) <= "00100000000111010000000000000000";
                        f_reg(348) <= "00010101011110010000000000100000";
                        f_reg(349) <= "10101111101010110000011101000100";
                        f_reg(350) <= "10001100000111010000011110010100";
                        f_reg(351) <= "00011111101000000000000000000011";
                        f_reg(352) <= "00100000000111010000000000111100";
                        f_reg(353) <= "00010000000000000000000000000010";
                        f_reg(354) <= "00100000000111010000000000000000";
                        f_reg(355) <= "00010101100110100000000000011001";
                        f_reg(356) <= "10101111101011000000011101001000";
                        f_reg(357) <= "10001100000111010000011110010100";
                        f_reg(358) <= "00011111101000000000000000000011";
                        f_reg(359) <= "00100000000111010000000000111100";
                        f_reg(360) <= "00010000000000000000000000000010";
                        f_reg(361) <= "00100000000111010000000000000000";
                        f_reg(362) <= "00010101101110110000000000010010";
                        f_reg(363) <= "10101111101011010000011101001100";
                        f_reg(364) <= "10001100000111010000011110010100";
                        f_reg(365) <= "00011111101000000000000000000011";
                        f_reg(366) <= "00100000000111010000000000111100";
                        f_reg(367) <= "00010000000000000000000000000010";
                        f_reg(368) <= "00100000000111010000000000000000";
                        f_reg(369) <= "00010101110111000000000000001011";
                        f_reg(370) <= "10101111101011100000011101010000";
                        f_reg(371) <= "10001100000111010000011110010100";
                        f_reg(372) <= "00011111101000000000000000000011";
                        f_reg(373) <= "00100000000111010000000000111100";
                        f_reg(374) <= "00010000000000000000000000000010";
                        f_reg(375) <= "00100000000111010000000000000000";
                        f_reg(376) <= "00010111110111110000000000000100";
                        f_reg(377) <= "10101111101111100000011101010100";
                        f_reg(378) <= "10101100000111010000011110010100";
                        f_reg(379) <= "00010000000000001111111110001000";
                        f_reg(380) <= "10001100000111010000011110010100";
                        f_reg(381) <= "10001111101000010000011100011100";
                        f_reg(382) <= "10001100000111010000011110010100";
                        f_reg(383) <= "10001111101011110000011100011100";
                        f_reg(384) <= "00010100001011111111111111111100";
                        f_reg(385) <= "10001100000111010000011110010100";
                        f_reg(386) <= "10001111101000100000011100100000";
                        f_reg(387) <= "10001100000111010000011110010100";
                        f_reg(388) <= "10001111101100000000011100100000";
                        f_reg(389) <= "00010100010100001111111111111100";
                        f_reg(390) <= "10001100000111010000011110010100";
                        f_reg(391) <= "10001111101000110000011100100100";
                        f_reg(392) <= "10001100000111010000011110010100";
                        f_reg(393) <= "10001111101100010000011100100100";
                        f_reg(394) <= "00010100011100011111111111111100";
                        f_reg(395) <= "10001100000111010000011110010100";
                        f_reg(396) <= "10001111101001000000011100101000";
                        f_reg(397) <= "10001100000111010000011110010100";
                        f_reg(398) <= "10001111101100100000011100101000";
                        f_reg(399) <= "00010100100100101111111111111100";
                        f_reg(400) <= "10001100000111010000011110010100";
                        f_reg(401) <= "10001111101001010000011100101100";
                        f_reg(402) <= "10001100000111010000011110010100";
                        f_reg(403) <= "10001111101100110000011100101100";
                        f_reg(404) <= "00010100101100111111111111111100";
                        f_reg(405) <= "10001100000111010000011110010100";
                        f_reg(406) <= "10001111101001100000011100110000";
                        f_reg(407) <= "10001100000111010000011110010100";
                        f_reg(408) <= "10001111101101000000011100110000";
                        f_reg(409) <= "00010100110101001111111111111100";
                        f_reg(410) <= "10001100000111010000011110010100";
                        f_reg(411) <= "10001111101001110000011100110100";
                        f_reg(412) <= "10001100000111010000011110010100";
                        f_reg(413) <= "10001111101101010000011100110100";
                        f_reg(414) <= "00010100111101011111111111111100";
                        f_reg(415) <= "10001100000111010000011110010100";
                        f_reg(416) <= "10001111101010000000011100111000";
                        f_reg(417) <= "10001100000111010000011110010100";
                        f_reg(418) <= "10001111101101100000011100111000";
                        f_reg(419) <= "00010101000101101111111111111100";
                        f_reg(420) <= "10001100000111010000011110010100";
                        f_reg(421) <= "10001111101010010000011100111100";
                        f_reg(422) <= "10001100000111010000011110010100";
                        f_reg(423) <= "10001111101101110000011100111100";
                        f_reg(424) <= "00010101001101111111111111111100";
                        f_reg(425) <= "10001100000111010000011110010100";
                        f_reg(426) <= "10001111101010100000011101000000";
                        f_reg(427) <= "10001100000111010000011110010100";
                        f_reg(428) <= "10001111101110000000011101000000";
                        f_reg(429) <= "00010101010110001111111111111100";
                        f_reg(430) <= "10001100000111010000011110010100";
                        f_reg(431) <= "10001111101010110000011101000100";
                        f_reg(432) <= "10001100000111010000011110010100";
                        f_reg(433) <= "10001111101110010000011101000100";
                        f_reg(434) <= "00010101011110011111111111111100";
                        f_reg(435) <= "10001100000111010000011110010100";
                        f_reg(436) <= "10001111101011000000011101001000";
                        f_reg(437) <= "10001100000111010000011110010100";
                        f_reg(438) <= "10001111101110100000011101001000";
                        f_reg(439) <= "00010101100110101111111111111100";
                        f_reg(440) <= "10001100000111010000011110010100";
                        f_reg(441) <= "10001111101011010000011101001100";
                        f_reg(442) <= "10001100000111010000011110010100";
                        f_reg(443) <= "10001111101110110000011101001100";
                        f_reg(444) <= "00010101101110111111111111111100";
                        f_reg(445) <= "10001100000111010000011110010100";
                        f_reg(446) <= "10001111101011100000011101010000";
                        f_reg(447) <= "10001100000111010000011110010100";
                        f_reg(448) <= "10001111101111000000011101010000";
                        f_reg(449) <= "00010101110111001111111111111100";
                        f_reg(450) <= "10001100000111010000011110010100";
                        f_reg(451) <= "10001111101111100000011101010100";
                        f_reg(452) <= "10001100000111010000011110010100";
                        f_reg(453) <= "10001111101111110000011101010100";
                        f_reg(454) <= "00010111110111111111111111111100";
                        f_reg(455) <= "00010000000000001111111100111100";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000001111100111";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011110001011000110";
                        f_reg(4) <= "00000000000000010001000000100011";
                        f_reg(5) <= "00110000010000110010110010110100";
                        f_reg(6) <= "00000000000000100010010111000011";
                        f_reg(7) <= "00000000100000110010100000100101";
                        f_reg(8) <= "00000000101001000011000000100111";
                        f_reg(9) <= "00000000000001000011100000100000";
                        f_reg(10) <= "00000000110001100100000000100110";
                        f_reg(11) <= "00000000011001110100100000000110";
                        f_reg(12) <= "00000000100001010101000000101011";
                        f_reg(13) <= "00111100000010111011000100000110";
                        f_reg(14) <= "00000000001000000110000000100111";
                        f_reg(15) <= "00000000000000000000000000000000";
                        f_reg(16) <= "00000000100010110110100000100001";
                        f_reg(17) <= "00000000100000100111000000100100";
                        f_reg(18) <= "00000001110010010111100000000111";
                        f_reg(19) <= "00000000000010101000010101000011";
                        f_reg(20) <= "00000001110010011000100000100110";
                        f_reg(21) <= "00000001010011011001000000100001";
                        f_reg(22) <= "00111100000100111111100001001000";
                        f_reg(23) <= "00110000100101000010101000100001";
                        f_reg(24) <= "00110010001101011110100101000110";
                        f_reg(25) <= "00000000000001000010010101000011";
                        f_reg(26) <= "00110001011101100000001011101110";
                        f_reg(27) <= "00000001111001111011100000100011";
                        f_reg(28) <= "00000000000000000000000000000000";
                        f_reg(29) <= "00000010000000111100000000100010";
                        f_reg(30) <= "00000010101101111100100000100101";
                        f_reg(31) <= "00000001110100101101000000100111";
                        f_reg(32) <= "00000000101011101101100000100101";
                        f_reg(33) <= "00000011001000111110000000000110";
                        f_reg(34) <= "00110011100111010110101000011011";
                        f_reg(35) <= "00000010101101111111000000100101";
                        f_reg(36) <= "00100011000001101011100111011001";
                        f_reg(37) <= "00000000000100110000110101000011";
                        f_reg(38) <= "00111100000000101011111011010101";
                        f_reg(39) <= "00000001011110110100100000100101";
                        f_reg(40) <= "00000011010000010101000000100000";
                        f_reg(41) <= "00000001010101000110100000100001";
                        f_reg(42) <= "00101101101100010110111101000101";
                        f_reg(43) <= "00000000110111010111100000000111";
                        f_reg(44) <= "00000010010011110011100000100100";
                        f_reg(45) <= "00000000010100011000000000100101";
                        f_reg(46) <= "00000010110100000010100000100110";
                        f_reg(47) <= "00101110110011100011000111001011";
                        f_reg(48) <= "00101001000000111100000010111011";
                        f_reg(49) <= "00000000101001101110000000100001";
                        f_reg(50) <= "00000011011011001010100000100110";
                        f_reg(51) <= "00000010101111101011100000101011";
                        f_reg(52) <= "00000000000000000000000000000000";
                        f_reg(53) <= "00000000111001001100000000000111";
                        f_reg(54) <= "10101100000010000000010000011100";
                        f_reg(55) <= "00000001011011101001100000100110";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000111101000111000010";
                        f_reg(58) <= "00000000000111000000111001000011";
                        f_reg(59) <= "00100110111010101001000110111000";
                        f_reg(60) <= "10101100000110010000010000100000";
                        f_reg(61) <= "00110100101101001111111000101001";
                        f_reg(62) <= "00100011010011010010111110011100";
                        f_reg(63) <= "00000001001101001110100000100001";
                        f_reg(64) <= "00000000000000000000000000000000";
                        f_reg(65) <= "00000011000000001001000000101011";
                        f_reg(66) <= "00000011101000010111100000100101";
                        f_reg(67) <= "00000000000000000000000000000000";
                        f_reg(68) <= "00000001010011110001000000100111";
                        f_reg(69) <= "10101100000011010000010000100100";
                        f_reg(70) <= "10101100000100100000010000101000";
                        f_reg(71) <= "10101100000100110000010000101100";
                        f_reg(72) <= "00000000000000000000000000000000";
                        f_reg(73) <= "10101100000000100000010000110000";
                        f_reg(74) <= "00100011111111111111111111111111";
                        f_reg(75) <= "00011111111000001111111110111000";
                        f_reg(76) <= "00010000000000000000000110111101";
                        f_reg(77) <= "00111100000111100000001111100111";
                        f_reg(78) <= "00111100000111110000001111100111";
                        f_reg(79) <= "00000000000111101111010000000010";
                        f_reg(80) <= "00000000000111111111110000000010";
                        f_reg(81) <= "00111100000000011110001011000110";
                        f_reg(82) <= "00111100000011111110001011000110";
                        f_reg(83) <= "00000000000000010001000000100011";
                        f_reg(84) <= "00000000000011111000000000100011";
                        f_reg(85) <= "00110000010000110010110010110100";
                        f_reg(86) <= "00110010000100010010110010110100";
                        f_reg(87) <= "00000000000000100010010111000011";
                        f_reg(88) <= "00000000000100001001010111000011";
                        f_reg(89) <= "00000000100000110010100000100101";
                        f_reg(90) <= "00000010010100011001100000100101";
                        f_reg(91) <= "00000000101001000011000000100111";
                        f_reg(92) <= "00000010011100101010000000100111";
                        f_reg(93) <= "00000000000001000011100000100000";
                        f_reg(94) <= "00000000000100101010100000100000";
                        f_reg(95) <= "00000000110001100100000000100110";
                        f_reg(96) <= "00000010100101001011000000100110";
                        f_reg(97) <= "00000000011001110100100000000110";
                        f_reg(98) <= "00000010001101011011100000000110";
                        f_reg(99) <= "00000000100001010101000000101011";
                        f_reg(100) <= "00000010010100111100000000101011";
                        f_reg(101) <= "00111100000010111011000100000110";
                        f_reg(102) <= "00111100000110011011000100000110";
                        f_reg(103) <= "00000000001000000110000000100111";
                        f_reg(104) <= "00000001111000001101000000100111";
                        f_reg(105) <= "00000000000000000000000000000000";
                        f_reg(106) <= "00000000000000000000000000000000";
                        f_reg(107) <= "00000000100010110110100000100001";
                        f_reg(108) <= "00000010010110011101100000100001";
                        f_reg(109) <= "00000000100000100111000000100100";
                        f_reg(110) <= "00000010010100001110000000100100";
                        f_reg(111) <= "00000001110010010011000000000111";
                        f_reg(112) <= "00000011100101111010000000000111";
                        f_reg(113) <= "00000000000010100000110101000011";
                        f_reg(114) <= "00000000000110000111110101000011";
                        f_reg(115) <= "00000001110010010001000000100110";
                        f_reg(116) <= "00000011100101111000000000100110";
                        f_reg(117) <= "00000001010011010100100000100001";
                        f_reg(118) <= "00000011000110111011100000100001";
                        f_reg(119) <= "00111100000010101111100001001000";
                        f_reg(120) <= "00111100000110001111100001001000";
                        f_reg(121) <= "00110000100011010010101000100001";
                        f_reg(122) <= "00110010010110110010101000100001";
                        f_reg(123) <= "00010101011110010000000100000001";
                        f_reg(124) <= "10101100000010110000010000110100";
                        f_reg(125) <= "00110000010010111110100101000110";
                        f_reg(126) <= "00110010000110011110100101000110";
                        f_reg(127) <= "00000000000001000010010101000011";
                        f_reg(128) <= "00000000000100101001010101000011";
                        f_reg(129) <= "10001100000000100000010000110100";
                        f_reg(130) <= "10001100000100000000010000110100";
                        f_reg(131) <= "00010100010100001111111111111110";
                        f_reg(132) <= "00010101000101100000000011111000";
                        f_reg(133) <= "10101100000010000000010000110100";
                        f_reg(134) <= "00110000010010000000001011101110";
                        f_reg(135) <= "00110010000101100000001011101110";
                        f_reg(136) <= "00010100010100000000000011110100";
                        f_reg(137) <= "10101100000000100000010000111000";
                        f_reg(138) <= "00000000110001110001000000100011";
                        f_reg(139) <= "00000010100101011000000000100011";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000000000000000000000000000";
                        f_reg(142) <= "00000000001000110011000000100010";
                        f_reg(143) <= "00000001111100011010000000100010";
                        f_reg(144) <= "00000001011000100011100000100101";
                        f_reg(145) <= "00000011001100001010100000100101";
                        f_reg(146) <= "00000001110010010000100000100111";
                        f_reg(147) <= "00000011100101110111100000100111";
                        f_reg(148) <= "00010100111101010000000011101000";
                        f_reg(149) <= "10101100000001110000010000111100";
                        f_reg(150) <= "00000000101011100011100000100101";
                        f_reg(151) <= "00000010011111001010100000100101";
                        f_reg(152) <= "10001100000001010000010000111100";
                        f_reg(153) <= "10001100000100110000010000111100";
                        f_reg(154) <= "00010100101100111111111111111110";
                        f_reg(155) <= "00000000101000110111000000000110";
                        f_reg(156) <= "00000010011100011110000000000110";
                        f_reg(157) <= "00110001110000110110101000011011";
                        f_reg(158) <= "00110011100100010110101000011011";
                        f_reg(159) <= "00000001011000100111000000100101";
                        f_reg(160) <= "00000011001100001110000000100101";
                        f_reg(161) <= "00100000110010111011100111011001";
                        f_reg(162) <= "00100010100110011011100111011001";
                        f_reg(163) <= "00000000000010100001010101000011";
                        f_reg(164) <= "00000000000110001000010101000011";
                        f_reg(165) <= "00111100000001101011111011010101";
                        f_reg(166) <= "00111100000101001011111011010101";
                        f_reg(167) <= "10001100000010100000010000111000";
                        f_reg(168) <= "10001100000110000000010000111000";
                        f_reg(169) <= "00010101010110001111111111111110";
                        f_reg(170) <= "00010100101100110000000011010010";
                        f_reg(171) <= "10101100000001010000010000111000";
                        f_reg(172) <= "00000001010001110010100000100101";
                        f_reg(173) <= "00000011000101011001100000100101";
                        f_reg(174) <= "00010100101100110000000011001110";
                        f_reg(175) <= "10101100000001010000010000111100";
                        f_reg(176) <= "00000000001000100010100000100000";
                        f_reg(177) <= "00000001111100001001100000100000";
                        f_reg(178) <= "00000000101011010000100000100001";
                        f_reg(179) <= "00000010011110110111100000100001";
                        f_reg(180) <= "00101100001000100110111101000101";
                        f_reg(181) <= "00101101111100000110111101000101";
                        f_reg(182) <= "00000001011000110010100000000111";
                        f_reg(183) <= "00000011001100011001100000000111";
                        f_reg(184) <= "00000001001001010110100000100100";
                        f_reg(185) <= "00000010111100111101100000100100";
                        f_reg(186) <= "00000000110000100000100000100101";
                        f_reg(187) <= "00000010100100000111100000100101";
                        f_reg(188) <= "00000001000000010001100000100110";
                        f_reg(189) <= "00000010110011111000100000100110";
                        f_reg(190) <= "00101101000010010011000111001011";
                        f_reg(191) <= "00101110110101110011000111001011";
                        f_reg(192) <= "10001100000001010000010000110100";
                        f_reg(193) <= "10001100000100110000010000110100";
                        f_reg(194) <= "00010100101100111111111111111110";
                        f_reg(195) <= "00101000101001101100000010111011";
                        f_reg(196) <= "00101010011101001100000010111011";
                        f_reg(197) <= "00000000011010110001000000100001";
                        f_reg(198) <= "00000010001110011000000000100001";
                        f_reg(199) <= "00000000111011000000100000100110";
                        f_reg(200) <= "00000010101110100111100000100110";
                        f_reg(201) <= "00000000001011100100000000101011";
                        f_reg(202) <= "00000001111111001011000000101011";
                        f_reg(203) <= "00000000000000000000000000000000";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000001101001000101100000000111";
                        f_reg(206) <= "00000011011100101100100000000111";
                        f_reg(207) <= "00010100101100110000000010101101";
                        f_reg(208) <= "10101100000001010000010000011100";
                        f_reg(209) <= "00000001010010010011100000100110";
                        f_reg(210) <= "00000011000101111010100000100110";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000001100110000111000010";
                        f_reg(214) <= "00000000000101001101000111000010";
                        f_reg(215) <= "00000000000000100000111001000011";
                        f_reg(216) <= "00000000000100000111111001000011";
                        f_reg(217) <= "00100101000011101001000110111000";
                        f_reg(218) <= "00100110110111001001000110111000";
                        f_reg(219) <= "10001100000001000000010000111000";
                        f_reg(220) <= "10001100000100100000010000111000";
                        f_reg(221) <= "00010100100100101111111111111110";
                        f_reg(222) <= "00010100100100100000000010011110";
                        f_reg(223) <= "10101100000001000000010000100000";
                        f_reg(224) <= "00110100011011011111111000101001";
                        f_reg(225) <= "00110110001110111111111000101001";
                        f_reg(226) <= "00100001100001010010111110011100";
                        f_reg(227) <= "00100011010100110010111110011100";
                        f_reg(228) <= "10001100000010100000010000111100";
                        f_reg(229) <= "10001100000110000000010000111100";
                        f_reg(230) <= "00010101010110001111111111111110";
                        f_reg(231) <= "00000001010011010100100000100001";
                        f_reg(232) <= "00000011000110111011100000100001";
                        f_reg(233) <= "00000000000000000000000000000000";
                        f_reg(234) <= "00000000000000000000000000000000";
                        f_reg(235) <= "00000001011000000011000000101011";
                        f_reg(236) <= "00000011001000001010000000101011";
                        f_reg(237) <= "00000001001000010001000000100101";
                        f_reg(238) <= "00000010111011111000000000100101";
                        f_reg(239) <= "00000000000000000000000000000000";
                        f_reg(240) <= "00000000000000000000000000000000";
                        f_reg(241) <= "00000001110000100100000000100111";
                        f_reg(242) <= "00000011100100001011000000100111";
                        f_reg(243) <= "00010100101100110000000010001001";
                        f_reg(244) <= "10101100000001010000010000100100";
                        f_reg(245) <= "00010100110101000000000010000111";
                        f_reg(246) <= "10101100000001100000010000101000";
                        f_reg(247) <= "00010100111101010000000010000101";
                        f_reg(248) <= "10101100000001110000010000101100";
                        f_reg(249) <= "00000000000000000000000000000000";
                        f_reg(250) <= "00000000000000000000000000000000";
                        f_reg(251) <= "00010101000101100000000010000001";
                        f_reg(252) <= "10101100000010000000010000110000";
                        f_reg(253) <= "00100011110111011111111100000110";
                        f_reg(254) <= "00010011101000000000000000010011";
                        f_reg(255) <= "00100011110111011111111000001100";
                        f_reg(256) <= "00010011101000000000000000010001";
                        f_reg(257) <= "00100011110111011111110100010010";
                        f_reg(258) <= "00010011101000000000000000001111";
                        f_reg(259) <= "00100011110111101111111111111111";
                        f_reg(260) <= "00100011111111111111111111111111";
                        f_reg(261) <= "00010111110111110000000001110111";
                        f_reg(262) <= "00011111111000001111111101001011";
                        f_reg(263) <= "00010000000000000000000100000010";
                        f_reg(264) <= "00000000000000000000000000000000";
                        f_reg(265) <= "00000000000000000000000000000000";
                        f_reg(266) <= "00000000000000000000000000000000";
                        f_reg(267) <= "00000000000000000000000000000000";
                        f_reg(268) <= "00000000000000000000000000000000";
                        f_reg(269) <= "00000000000000000000000000000000";
                        f_reg(270) <= "00000000000000000000000000000000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "10001100000111010000011110010100";
                        f_reg(274) <= "00011111101000000000000000000011";
                        f_reg(275) <= "00100000000111010000000000111100";
                        f_reg(276) <= "00010000000000000000000000000010";
                        f_reg(277) <= "00100000000111010000000000000000";
                        f_reg(278) <= "00010100001011110000000001100110";
                        f_reg(279) <= "10101111101000010000011100011100";
                        f_reg(280) <= "10001100000111010000011110010100";
                        f_reg(281) <= "00011111101000000000000000000011";
                        f_reg(282) <= "00100000000111010000000000111100";
                        f_reg(283) <= "00010000000000000000000000000010";
                        f_reg(284) <= "00100000000111010000000000000000";
                        f_reg(285) <= "00010100010100000000000001011111";
                        f_reg(286) <= "10101111101000100000011100100000";
                        f_reg(287) <= "10001100000111010000011110010100";
                        f_reg(288) <= "00011111101000000000000000000011";
                        f_reg(289) <= "00100000000111010000000000111100";
                        f_reg(290) <= "00010000000000000000000000000010";
                        f_reg(291) <= "00100000000111010000000000000000";
                        f_reg(292) <= "00010100011100010000000001011000";
                        f_reg(293) <= "10101111101000110000011100100100";
                        f_reg(294) <= "10001100000111010000011110010100";
                        f_reg(295) <= "00011111101000000000000000000011";
                        f_reg(296) <= "00100000000111010000000000111100";
                        f_reg(297) <= "00010000000000000000000000000010";
                        f_reg(298) <= "00100000000111010000000000000000";
                        f_reg(299) <= "00010100100100100000000001010001";
                        f_reg(300) <= "10101111101001000000011100101000";
                        f_reg(301) <= "10001100000111010000011110010100";
                        f_reg(302) <= "00011111101000000000000000000011";
                        f_reg(303) <= "00100000000111010000000000111100";
                        f_reg(304) <= "00010000000000000000000000000010";
                        f_reg(305) <= "00100000000111010000000000000000";
                        f_reg(306) <= "00010100101100110000000001001010";
                        f_reg(307) <= "10101111101001010000011100101100";
                        f_reg(308) <= "10001100000111010000011110010100";
                        f_reg(309) <= "00011111101000000000000000000011";
                        f_reg(310) <= "00100000000111010000000000111100";
                        f_reg(311) <= "00010000000000000000000000000010";
                        f_reg(312) <= "00100000000111010000000000000000";
                        f_reg(313) <= "00010100110101000000000001000011";
                        f_reg(314) <= "10101111101001100000011100110000";
                        f_reg(315) <= "10001100000111010000011110010100";
                        f_reg(316) <= "00011111101000000000000000000011";
                        f_reg(317) <= "00100000000111010000000000111100";
                        f_reg(318) <= "00010000000000000000000000000010";
                        f_reg(319) <= "00100000000111010000000000000000";
                        f_reg(320) <= "00010100111101010000000000111100";
                        f_reg(321) <= "10101111101001110000011100110100";
                        f_reg(322) <= "10001100000111010000011110010100";
                        f_reg(323) <= "00011111101000000000000000000011";
                        f_reg(324) <= "00100000000111010000000000111100";
                        f_reg(325) <= "00010000000000000000000000000010";
                        f_reg(326) <= "00100000000111010000000000000000";
                        f_reg(327) <= "00010101000101100000000000110101";
                        f_reg(328) <= "10101111101010000000011100111000";
                        f_reg(329) <= "10001100000111010000011110010100";
                        f_reg(330) <= "00011111101000000000000000000011";
                        f_reg(331) <= "00100000000111010000000000111100";
                        f_reg(332) <= "00010000000000000000000000000010";
                        f_reg(333) <= "00100000000111010000000000000000";
                        f_reg(334) <= "00010101001101110000000000101110";
                        f_reg(335) <= "10101111101010010000011100111100";
                        f_reg(336) <= "10001100000111010000011110010100";
                        f_reg(337) <= "00011111101000000000000000000011";
                        f_reg(338) <= "00100000000111010000000000111100";
                        f_reg(339) <= "00010000000000000000000000000010";
                        f_reg(340) <= "00100000000111010000000000000000";
                        f_reg(341) <= "00010101010110000000000000100111";
                        f_reg(342) <= "10101111101010100000011101000000";
                        f_reg(343) <= "10001100000111010000011110010100";
                        f_reg(344) <= "00011111101000000000000000000011";
                        f_reg(345) <= "00100000000111010000000000111100";
                        f_reg(346) <= "00010000000000000000000000000010";
                        f_reg(347) <= "00100000000111010000000000000000";
                        f_reg(348) <= "00010101011110010000000000100000";
                        f_reg(349) <= "10101111101010110000011101000100";
                        f_reg(350) <= "10001100000111010000011110010100";
                        f_reg(351) <= "00011111101000000000000000000011";
                        f_reg(352) <= "00100000000111010000000000111100";
                        f_reg(353) <= "00010000000000000000000000000010";
                        f_reg(354) <= "00100000000111010000000000000000";
                        f_reg(355) <= "00010101100110100000000000011001";
                        f_reg(356) <= "10101111101011000000011101001000";
                        f_reg(357) <= "10001100000111010000011110010100";
                        f_reg(358) <= "00011111101000000000000000000011";
                        f_reg(359) <= "00100000000111010000000000111100";
                        f_reg(360) <= "00010000000000000000000000000010";
                        f_reg(361) <= "00100000000111010000000000000000";
                        f_reg(362) <= "00010101101110110000000000010010";
                        f_reg(363) <= "10101111101011010000011101001100";
                        f_reg(364) <= "10001100000111010000011110010100";
                        f_reg(365) <= "00011111101000000000000000000011";
                        f_reg(366) <= "00100000000111010000000000111100";
                        f_reg(367) <= "00010000000000000000000000000010";
                        f_reg(368) <= "00100000000111010000000000000000";
                        f_reg(369) <= "00010101110111000000000000001011";
                        f_reg(370) <= "10101111101011100000011101010000";
                        f_reg(371) <= "10001100000111010000011110010100";
                        f_reg(372) <= "00011111101000000000000000000011";
                        f_reg(373) <= "00100000000111010000000000111100";
                        f_reg(374) <= "00010000000000000000000000000010";
                        f_reg(375) <= "00100000000111010000000000000000";
                        f_reg(376) <= "00010111110111110000000000000100";
                        f_reg(377) <= "10101111101111100000011101010100";
                        f_reg(378) <= "10101100000111010000011110010100";
                        f_reg(379) <= "00010000000000001111111110001000";
                        f_reg(380) <= "10001100000111010000011110010100";
                        f_reg(381) <= "10001111101000010000011100011100";
                        f_reg(382) <= "10001100000111010000011110010100";
                        f_reg(383) <= "10001111101011110000011100011100";
                        f_reg(384) <= "00010100001011111111111111111100";
                        f_reg(385) <= "10001100000111010000011110010100";
                        f_reg(386) <= "10001111101000100000011100100000";
                        f_reg(387) <= "10001100000111010000011110010100";
                        f_reg(388) <= "10001111101100000000011100100000";
                        f_reg(389) <= "00010100010100001111111111111100";
                        f_reg(390) <= "10001100000111010000011110010100";
                        f_reg(391) <= "10001111101000110000011100100100";
                        f_reg(392) <= "10001100000111010000011110010100";
                        f_reg(393) <= "10001111101100010000011100100100";
                        f_reg(394) <= "00010100011100011111111111111100";
                        f_reg(395) <= "10001100000111010000011110010100";
                        f_reg(396) <= "10001111101001000000011100101000";
                        f_reg(397) <= "10001100000111010000011110010100";
                        f_reg(398) <= "10001111101100100000011100101000";
                        f_reg(399) <= "00010100100100101111111111111100";
                        f_reg(400) <= "10001100000111010000011110010100";
                        f_reg(401) <= "10001111101001010000011100101100";
                        f_reg(402) <= "10001100000111010000011110010100";
                        f_reg(403) <= "10001111101100110000011100101100";
                        f_reg(404) <= "00010100101100111111111111111100";
                        f_reg(405) <= "10001100000111010000011110010100";
                        f_reg(406) <= "10001111101001100000011100110000";
                        f_reg(407) <= "10001100000111010000011110010100";
                        f_reg(408) <= "10001111101101000000011100110000";
                        f_reg(409) <= "00010100110101001111111111111100";
                        f_reg(410) <= "10001100000111010000011110010100";
                        f_reg(411) <= "10001111101001110000011100110100";
                        f_reg(412) <= "10001100000111010000011110010100";
                        f_reg(413) <= "10001111101101010000011100110100";
                        f_reg(414) <= "00010100111101011111111111111100";
                        f_reg(415) <= "10001100000111010000011110010100";
                        f_reg(416) <= "10001111101010000000011100111000";
                        f_reg(417) <= "10001100000111010000011110010100";
                        f_reg(418) <= "10001111101101100000011100111000";
                        f_reg(419) <= "00010101000101101111111111111100";
                        f_reg(420) <= "10001100000111010000011110010100";
                        f_reg(421) <= "10001111101010010000011100111100";
                        f_reg(422) <= "10001100000111010000011110010100";
                        f_reg(423) <= "10001111101101110000011100111100";
                        f_reg(424) <= "00010101001101111111111111111100";
                        f_reg(425) <= "10001100000111010000011110010100";
                        f_reg(426) <= "10001111101010100000011101000000";
                        f_reg(427) <= "10001100000111010000011110010100";
                        f_reg(428) <= "10001111101110000000011101000000";
                        f_reg(429) <= "00010101010110001111111111111100";
                        f_reg(430) <= "10001100000111010000011110010100";
                        f_reg(431) <= "10001111101010110000011101000100";
                        f_reg(432) <= "10001100000111010000011110010100";
                        f_reg(433) <= "10001111101110010000011101000100";
                        f_reg(434) <= "00010101011110011111111111111100";
                        f_reg(435) <= "10001100000111010000011110010100";
                        f_reg(436) <= "10001111101011000000011101001000";
                        f_reg(437) <= "10001100000111010000011110010100";
                        f_reg(438) <= "10001111101110100000011101001000";
                        f_reg(439) <= "00010101100110101111111111111100";
                        f_reg(440) <= "10001100000111010000011110010100";
                        f_reg(441) <= "10001111101011010000011101001100";
                        f_reg(442) <= "10001100000111010000011110010100";
                        f_reg(443) <= "10001111101110110000011101001100";
                        f_reg(444) <= "00010101101110111111111111111100";
                        f_reg(445) <= "10001100000111010000011110010100";
                        f_reg(446) <= "10001111101011100000011101010000";
                        f_reg(447) <= "10001100000111010000011110010100";
                        f_reg(448) <= "10001111101111000000011101010000";
                        f_reg(449) <= "00010101110111001111111111111100";
                        f_reg(450) <= "10001100000111010000011110010100";
                        f_reg(451) <= "10001111101111100000011101010100";
                        f_reg(452) <= "10001100000111010000011110010100";
                        f_reg(453) <= "10001111101111110000011101010100";
                        f_reg(454) <= "00010111110111111111111111111100";
                        f_reg(455) <= "00010000000000001111111100111100";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                        f_reg(466) <= "00000000000000000000000000000000";
                        f_reg(467) <= "00000000000000000000000000000000";
                        f_reg(468) <= "00000000000000000000000000000000";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000001111100111";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test59_Reg_COMBINED;
