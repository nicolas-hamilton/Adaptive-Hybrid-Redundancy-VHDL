--| Comparator_TB.vhd
--| Test the functionality of the comparator
library IEEE;
use IEEE.std_logic_1164.all;

entity Comparator_TB is
end Comparator_TB;

architecture testbench of Comparator_TB is
--| Declare Components
	component Comparator is
		port (i_S			: in  std_logic_vector(31 downto 0);
				i_NAND_AB		: in  std_logic;
				i_OR_AB		: in  std_logic;
				i_XNOR_AB		: in  std_logic;
				i_unsigned	: in  std_logic;
				i_COMP_SEL	: in  std_logic_vector(2 downto 0);
				o_Z			: out std_logic);
	end component;
	
	--| Declare Signals
	signal w_S : std_logic_vector(31 downto 0) := (others => '0');
	signal w_A : std_logic := '0';
	signal w_B : std_logic := '0';
	signal w_NAND_AB : std_logic;
	signal w_OR_AB : std_logic;
	signal w_XNOR_AB : std_logic;
	signal w_unsigned : std_logic := '0';
	signal w_COMP_SEL : std_logic_vector(2 downto 0) := (others => '0');
	signal w_Z : std_logic;
begin
	w_NAND_AB <= w_A NAND w_B;
	w_OR_AB <= w_A OR w_B;
	w_XNOR_AB <= w_A XNOR w_B;
	u_Comparator: Comparator
	port map (i_S => w_S,
				 i_NAND_AB => w_NAND_AB,
				 i_OR_AB => w_OR_AB,
				 i_XNOR_AB => w_XNOR_AB,
				 i_unsigned => w_UNSIGNED,
				 i_COMP_SEL => w_COMP_SEL,
				 o_Z => w_Z);
				 
	stimulus: process is
	begin
		-- Check all outputs for A=B=0, unsigned = 0
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=1, B=0, unsigned = 0
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=0, B=1, unsigned = 0
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '0';
		w_B <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=1, B=1, unsigned = 0
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=B=0, unsigned = 1
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '0';
		w_B <= '0';
		w_unsigned <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=1, B=0, unsigned = 1
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=0, B=1, unsigned = 1
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '0';
		w_B <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		
		-- Check all outputs for A=1, B=1, unsigned = 1
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= (others => '0');
		w_A <= '1';
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"0000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait for 20 ns;
		w_COMP_SEL <= B"000";
		w_S <= B"1000_0110_1000_0100_0001_0010_0100_0000";
		wait for 20 ns;
		w_COMP_SEL <= B"001";
		wait for 20 ns;
		w_COMP_SEL <= B"010";
		wait for 20 ns;
		w_COMP_SEL <= B"011";
		wait for 20 ns;
		w_COMP_SEL <= B"100";
		wait for 20 ns;
		w_COMP_SEL <= B"101";
		wait for 20 ns;
		w_COMP_SEL <= B"110";
		wait for 20 ns;
		w_COMP_SEL <= B"111";
		wait;
	end process stimulus;
end testbench;