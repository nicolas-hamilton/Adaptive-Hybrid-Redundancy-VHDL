--| Instruction_Dec_Enc.vhd
--| Decodes the 32-bit MIPS instruction to determine which portions of the ALU to activate.
--| Encodes some of these signals to control muxes in the datapath.
--|
--| INPUTS:
--| i_instr31 			- Instruction inputs
--| ...
--| i_instr00 			- Instruction inputs
--| i_BRANCH_OVERRIDE- Modify ALU_SRC_A(1) so that the ALU will use the PC input for ALU_SRC_A.
--|						- Override ALU_SRC_B and ALU_INV_B controls generated by decoding the
--|						  instruction.  Used by the controller to modify the behavior of the
--|						  datapath during the second cycle of a branch instruction.
--|						- Modify ALU_OUTPUT to select the adder output.  Used in the second cycle
--|						  of branch instructions to add the PC and the branch offset or 4.
--| i_DO_NOT_STORE	- Override the REG_SEL control generated by decoding the instruction.
--|						  Used by the controller to ensure data is only written to registers
--|						  during the write phase of the particular instruction when the ALU
--|						  result or data from memory is ready to be sampled and stored.
--| i_PC_STORE			- Override the REG_SEL control generated by decoding the instruction.
--|						  Cause the output of the datapath to be stored to the PC register.
--|						  Used for branch instructions to store the result of a branch to
--|						  the PC register.
--|						
--|
--| OUTPUTS:
--| o_ALU_SRC_A	- ALU Source A selector
--| o_ALU_SRC_B	- ALU Source B selector
--| o_ALU_INV_B	- ALU Invert B selector
--| o_COMP_SEL 	- Select the value to output from the Comparator
--| o_OVER_CTRL	- Select which overflow detection means should be used
--|					  (i.e. ADD, ADDI, SUB, or no overflow detection).
--| o_ALU_OUTPUT	- Select which ALU function should be output
--|						0 - Shift Left
--|						1 - Shift Right
--|						2 - Adder
--|						3 - AND
--|						4 - OR
--|						5 - XOR
--|						6 - NOR
--|						7 - Comparator
--|						8 - LUI
--|						9, 10, 11, 12, 13, 14, 15 - Shift Left
--| o_REG_SEL		- Select the destination register.
--| o_UNSIGNED		- Determine if the comparator is comparing sigend numbers (0) or unsigned
--|					  numbers (1).
--| o_overflow		- Determine if the comparator is performing a Less Than comparison that will
--|                 or will not produce an overflow.  No overflow can occur in BLTZ instructions,
--|					  but overflow can occur in SLT, SLTU, SLTI, and SLTIU instructions.  0 - no
--|					  overflow can occur, 1 - overflow can occur
--| o_imm_extend		- Determine if the immediate value should be 0 extended or sign extended
--| o_FSM_CTRL		- Finite State Machine Control Signal
--| o_INVALID_INSTR	- Signals when an invalid instruction is received
library IEEE;
use IEEE.std_logic_1164.all;

entity Instruction_Dec_Enc is
	port (i_instr31			: in  std_logic;
			i_instr30			: in  std_logic;
			i_instr29			: in  std_logic;
			i_instr28			: in  std_logic;
			i_instr27			: in  std_logic;
			i_instr26			: in  std_logic;
			i_instr20			: in  std_logic;
			i_instr19			: in  std_logic;
			i_instr18			: in  std_logic;
			i_instr17			: in  std_logic;
			i_instr16			: in  std_logic;
			i_instr05			: in  std_logic;
			i_instr04			: in  std_logic;
			i_instr03			: in  std_logic;
			i_instr02			: in  std_logic;
			i_instr01			: in  std_logic;
			i_instr00			: in  std_logic;
			i_BRANCH_OVERRIDE	: in  std_logic;
			i_DO_NOT_STORE		: in  std_logic;
			i_PC_STORE			: in  std_logic;
			o_ALU_SRC_A			: out std_logic_vector(1 downto 0);
			o_ALU_SRC_B			: out std_logic_vector(1 downto 0);
			o_ALU_INV_B 		: out std_logic;
			o_COMP_SEL			: out std_logic_vector(2 downto 0);
			o_OVER_CTRL 		: out std_logic_vector(1 downto 0);
			o_ALU_OUTPUT		: out std_logic_vector(3 downto 0);
			o_REG_SEL			: out std_logic_vector(1 downto 0);
			o_UNSIGNED			: out std_logic;
			o_overflow			: out std_logic;
			o_imm_extend		: out std_logic;
			o_FSM_CTRL			: out std_logic_vector(1 downto 0);
			o_INVALID_INSTR	: out std_logic);
end Instruction_Dec_Enc;

architecture a_Instruction_Dec_Enc of Instruction_Dec_Enc is
--| Define Components
	component myMUX2_N is
		generic (m_width : integer := 2);
		port (i_0 : in  std_logic_vector(m_width-1 downto 0);
				i_1 : in  std_logic_vector(m_width-1 downto 0);
				i_S : in  std_logic;
				o_Z : out std_logic_vector(m_width-1 downto 0));
	end component;
	
	component myMUX2_1 is
		port (i_0 : in  std_logic;
				i_1 : in  std_logic;
				i_S : in  std_logic;
				o_Z : out std_logic);
	end component;
	
	component Instruction_Decoder is
		port (i_instr31		: in  std_logic;
				i_instr30		: in  std_logic;
				i_instr29		: in  std_logic;
				i_instr28		: in  std_logic;
				i_instr27		: in  std_logic;
				i_instr26		: in  std_logic;
				i_instr20		: in  std_logic;
				i_instr19		: in  std_logic;
				i_instr18		: in  std_logic;
				i_instr17		: in  std_logic;
				i_instr16		: in  std_logic;
				i_instr05		: in  std_logic;
				i_instr04		: in  std_logic;
				i_instr03		: in  std_logic;
				i_instr02		: in  std_logic;
				i_instr01		: in  std_logic;
				i_instr00		: in  std_logic;
				o_ALU_SRC_A0	: out std_logic;
				o_ALU_SRC_B		: out std_logic_vector(1 downto 0);
				o_INV_B			: out std_logic;
				o_LTZ				: out std_logic;
				o_EQ				: out std_logic;
				o_NE				: out std_logic;
				o_LEZ				: out std_logic;
				o_GTZ				: out std_logic;
				o_RIGHT_SHIFT	: out std_logic;
				o_ADDER			: out std_logic;
				o_AND				: out std_logic;
				o_OR				: out std_logic;
				o_XOR				: out std_logic;
				o_NOR				: out std_logic;
				o_COMPARE		: out std_logic;
				o_LUI				: out std_logic;
				o_REG_SEL		: out std_logic_vector(1 downto 0);
				o_OVER_CTRL		: out std_logic_vector(1 downto 0);
				o_UNSIGNED		: out std_logic;
				o_overflow		: out std_logic;
				o_imm_extend	: out std_logic;
				o_FSM_CTRL		: out std_logic_vector(1 downto 0);
				o_INVALID_INSTR: out std_logic);
	end component;
	
	component Encoder6_3 is
		port (i_1 : in  std_logic;
				i_2 : in  std_logic;
				i_3 : in  std_logic;
				i_4 : in  std_logic;
				i_5 : in  std_logic;
				o_Z : out std_logic_vector(2 downto 0));
	end component;
	
	component Encoder9_4 is
		port (i_1 : in  std_logic;
				i_2 : in  std_logic;
				i_3 : in  std_logic;
				i_4 : in  std_logic;
				i_5 : in  std_logic;
				i_6 : in  std_logic;
				i_7 : in  std_logic;
				i_8 : in  std_logic;
				o_Z : out std_logic_vector(3 downto 0));
	end component;

--| Define Signals
	signal w_ALU_SRC_B	: std_logic_vector(1 downto 0);
	signal w_ALU_INV_B			: std_logic;
	signal w_LTZ			: std_logic;
	signal w_EQ				: std_logic;
	signal w_NE				: std_logic;
	signal w_LEZ			: std_logic;
	signal w_GTZ			: std_logic;
	signal w_RIGHT_SHIFT	: std_logic;
	signal w_ADDER			: std_logic;
	signal w_AND			: std_logic;
	signal w_OR				: std_logic;
	signal w_XOR			: std_logic;
	signal w_NOR			: std_logic;
	signal w_COMPARE		: std_logic;
	signal w_LUI			: std_logic;
	signal w_REG_SEL0, w_REG_SEL1		: std_logic_vector(1 downto 0);
	signal w_ALU_OUTPUT	: std_logic_vector(3 downto 0);
	
--| Define Constants
	constant k_one2 : std_logic_vector(1 downto 0) := B"11";
	constant k_zero1 : std_logic := '0';
	constant k_zero2 : std_logic_vector(1 downto 0) := B"00";
	constant k_two4 : std_logic_vector(3 downto 0) := B"0010";
	
begin
	o_ALU_SRC_A(1) <= i_BRANCH_OVERRIDE;
	
	-- Connect the Instruction Decoder
	u_Instruction_Decoder: Instruction_Decoder
	port map (i_instr31 => i_instr31,
				 i_instr30 => i_instr30,
				 i_instr29 => i_instr29,
				 i_instr28 => i_instr28,
				 i_instr27 => i_instr27,
				 i_instr26 => i_instr26,
				 i_instr20 => i_instr20,
				 i_instr19 => i_instr19,
				 i_instr18 => i_instr18,
				 i_instr17 => i_instr17,
				 i_instr16 => i_instr16,
				 i_instr05 => i_instr05,
				 i_instr04 => i_instr04,
				 i_instr03 => i_instr03,
				 i_instr02 => i_instr02,
				 i_instr01 => i_instr01,
				 i_instr00 => i_instr00,
				 o_ALU_SRC_A0 => o_ALU_SRC_A(0),
				 o_ALU_SRC_B => w_ALU_SRC_B,
				 o_INV_B => w_ALU_INV_B,
				 o_LTZ => w_LTZ,
				 o_EQ => w_EQ,
				 o_NE => w_NE,
				 o_LEZ => w_LEZ,
				 o_GTZ => w_GTZ,
				 o_RIGHT_SHIFT => w_RIGHT_SHIFT,
				 o_ADDER => w_ADDER,
				 o_AND => w_AND,
				 o_OR => w_OR,
				 o_XOR => w_XOR,
				 o_NOR => w_NOR,
				 o_COMPARE => w_COMPARE,
				 o_LUI => w_LUI,
				 o_REG_SEL => w_REG_SEL0,
				 o_OVER_CTRL => o_OVER_CTRL,
				 o_UNSIGNED => o_UNSIGNED,
				 o_overflow => o_overflow,
				 o_imm_extend => o_imm_extend,
				 o_FSM_CTRL => o_FSM_CTRL,
				 o_INVALID_INSTR => o_INVALID_INSTR);
		
	-- Encode the COMP_SEL signal
	u_Encoder6_3 : Encoder6_3
	port map (
		i_1 => w_LTZ,
		i_2 => w_EQ,
		i_3 => w_NE,
		i_4 => w_LEZ,
		i_5 => w_GTZ,
		o_Z => o_COMP_SEL);
		
	-- Encode the ALU_OUTPUT signal
	u_Encoder9_4 : Encoder9_4
	port map (
		i_1 => w_RIGHT_SHIFT,
		i_2 => w_ADDER,
		i_3 => w_AND,
		i_4 => w_OR,
		i_5 => w_XOR,
		i_6 => w_NOR,
		i_7 => w_COMPARE,
		i_8 => w_LUI,
		o_Z => w_ALU_OUTPUT);
	
	-- Determine whether ALU_SRC_B is dependent on the instruction or the current state
	u_myMUX2_SRC_B: myMUX2_N
	generic map (m_width => 2)
	port map (i_0 => w_ALU_SRC_B,
				 i_1 => k_one2,
				 i_S => i_BRANCH_OVERRIDE,
				 o_Z => o_ALU_SRC_B);
				 
	-- Determine whether ALU_INV_B is dependent on the instruction or the current state
	u_myMUX2_INV_B: myMUX2_1
	port map (i_0 => w_ALU_INV_B,
				 i_1 => k_zero1,
				 i_S => i_BRANCH_OVERRIDE,
				 o_Z => o_ALU_INV_B);
	
	-- Determine whether data should be written to the PC register
	u_myMUX2_REG_SEL1: myMUX2_N
	generic map (m_width => 2)
	port map (i_0 => w_REG_SEL0,
				 i_1 => k_one2,
				 i_S => i_PC_STORE,
				 o_Z => w_REG_SEL1);
				 
	-- Determine whether ALU_OUTPUT is dependent on the instruction or the current state
	u_myMUX2_ALU_OUTPUT: myMUX2_N
	generic map (m_width => 4)
	port map (i_0 => w_ALU_OUTPUT,
				 i_1 => k_two4,
				 i_S => i_BRANCH_OVERRIDE,
				 o_Z => o_ALU_OUTPUT);
	
	-- Determine whether data should be written to registers
	u_myMUX2_REG_SEL: myMUX2_N
	generic map (m_width => 2)
	port map (i_0 => w_REG_SEL1,
				 i_1 => k_zero2,
				 i_S => i_DO_NOT_STORE,
				 o_Z => o_REG_SEL);
	
end a_Instruction_Dec_Enc;