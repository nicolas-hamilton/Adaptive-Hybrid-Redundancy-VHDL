--| RIGHT_SHIFT.vhd
--| Implements the right shift function.  Shifts input A by the amount specified by SA.
--| Performs a logical right shift if w_fill is 0 and an arithmetic right shift if w_fill is 1.
--|
--| INPUTS:
--| i_A - Data Input
--| i_SA - Shift Amount
--| i_ARITH - 0 for logical shift, 1 for arithmetic shift
--|
--| OUTPUTS:
--| o_Z - Shifted input data (o_Z = i_A >> i_SA)
library IEEE;
use IEEE.std_logic_1164.all;

entity RIGHT_SHIFT is
	port (i_A		: in  std_logic_vector(31 downto 0);
			i_SA		: in  std_logic_vector(4 downto 0);
			i_ARITH	: in std_logic;
			o_Z		: out std_logic_vector(31 downto 0));
end RIGHT_SHIFT;

architecture a_RIGHT_SHIFT of RIGHT_SHIFT is
	-- Declare Components
	component myMUX2_1 is
		port (i_0 : in  std_logic;
				i_1 : in  std_logic;
				i_S : in  std_logic;
				o_Z : out std_logic
				);
	end component;
	
	component myMUX32_1 is
		port (i_0	: in  std_logic;
				i_1	: in  std_logic;
				i_2	: in  std_logic;
				i_3	: in  std_logic;
				i_4	: in  std_logic;
				i_5	: in  std_logic;
				i_6	: in  std_logic;
				i_7	: in  std_logic;
				i_8	: in  std_logic;
				i_9	: in  std_logic;
				i_10	: in  std_logic;
				i_11	: in  std_logic;
				i_12	: in  std_logic;
				i_13	: in  std_logic;
				i_14	: in  std_logic;
				i_15	: in  std_logic;
				i_16	: in  std_logic;
				i_17	: in  std_logic;
				i_18	: in  std_logic;
				i_19	: in  std_logic;
				i_20	: in  std_logic;
				i_21	: in  std_logic;
				i_22	: in  std_logic;
				i_23	: in  std_logic;
				i_24	: in  std_logic;
				i_25	: in  std_logic;
				i_26	: in  std_logic;
				i_27	: in  std_logic;
				i_28	: in  std_logic;
				i_29	: in  std_logic;
				i_30	: in  std_logic;
				i_31	: in  std_logic;
				i_S	: in  std_logic_vector (4 downto 0);
				o_Z	: out std_logic
				);
	end component;
	
	signal w_fill : std_logic;
	constant k_zero : std_logic := '0';

begin

	u_mux2_1 : myMUX2_1
	port map (i_0 => k_zero,
				 i_1 => i_A(31),
				 i_S => i_ARITH,
				 o_Z => w_fill);
	
	u_myMUX_bit31: myMUX32_1
	port map (i_0 => i_A(31),
				 i_1 => w_fill,
				 i_2 => w_fill,
				 i_3 => w_fill,
				 i_4 => w_fill,
				 i_5 => w_fill,
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(31));
	
	u_myMUX_bit30: myMUX32_1
	port map (i_0 => i_A(30),
				 i_1 => i_A(31),
				 i_2 => w_fill,
				 i_3 => w_fill,
				 i_4 => w_fill,
				 i_5 => w_fill,
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(30));
	
	u_myMUX_bit29: myMUX32_1
	port map (i_0 => i_A(29),
				 i_1 => i_A(30),
				 i_2 => i_A(31),
				 i_3 => w_fill,
				 i_4 => w_fill,
				 i_5 => w_fill,
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(29));
	
	u_myMUX_bit28: myMUX32_1
	port map (i_0 => i_A(28),
				 i_1 => i_A(29),
				 i_2 => i_A(30),
				 i_3 => i_A(31),
				 i_4 => w_fill,
				 i_5 => w_fill,
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(28));
	
	u_myMUX_bit27: myMUX32_1
	port map (i_0 => i_A(27),
				 i_1 => i_A(28),
				 i_2 => i_A(29),
				 i_3 => i_A(30),
				 i_4 => i_A(31),
				 i_5 => w_fill,
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(27));
	
	u_myMUX_bit26: myMUX32_1
	port map (i_0 => i_A(26),
				 i_1 => i_A(27),
				 i_2 => i_A(28),
				 i_3 => i_A(29),
				 i_4 => i_A(30),
				 i_5 => i_A(31),
				 i_6 => w_fill,
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(26));
	
	u_myMUX_bit25: myMUX32_1
	port map (i_0 => i_A(25),
				 i_1 => i_A(26),
				 i_2 => i_A(27),
				 i_3 => i_A(28),
				 i_4 => i_A(29),
				 i_5 => i_A(30),
				 i_6 => i_A(31),
				 i_7 => w_fill,
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(25));
	
	u_myMUX_bit24: myMUX32_1
	port map (i_0 => i_A(24),
				 i_1 => i_A(25),
				 i_2 => i_A(26),
				 i_3 => i_A(27),
				 i_4 => i_A(28),
				 i_5 => i_A(29),
				 i_6 => i_A(30),
				 i_7 => i_A(31),
				 i_8 => w_fill,
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(24));
	
	u_myMUX_bit23: myMUX32_1
	port map (i_0 => i_A(23),
				 i_1 => i_A(24),
				 i_2 => i_A(25),
				 i_3 => i_A(26),
				 i_4 => i_A(27),
				 i_5 => i_A(28),
				 i_6 => i_A(29),
				 i_7 => i_A(30),
				 i_8 => i_A(31),
				 i_9 => w_fill,
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(23));
	
	u_myMUX_bit22: myMUX32_1
	port map (i_0 => i_A(22),
				 i_1 => i_A(23),
				 i_2 => i_A(24),
				 i_3 => i_A(25),
				 i_4 => i_A(26),
				 i_5 => i_A(27),
				 i_6 => i_A(28),
				 i_7 => i_A(29),
				 i_8 => i_A(30),
				 i_9 => i_A(31),
				 i_10 => w_fill,
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(22));
	
	u_myMUX_bit21: myMUX32_1
	port map (i_0 => i_A(21),
				 i_1 => i_A(22),
				 i_2 => i_A(23),
				 i_3 => i_A(24),
				 i_4 => i_A(25),
				 i_5 => i_A(26),
				 i_6 => i_A(27),
				 i_7 => i_A(28),
				 i_8 => i_A(29),
				 i_9 => i_A(30),
				 i_10 => i_A(31),
				 i_11 => w_fill,
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(21));
	
	u_myMUX_bit20: myMUX32_1
	port map (i_0 => i_A(20),
				 i_1 => i_A(21),
				 i_2 => i_A(22),
				 i_3 => i_A(23),
				 i_4 => i_A(24),
				 i_5 => i_A(25),
				 i_6 => i_A(26),
				 i_7 => i_A(27),
				 i_8 => i_A(28),
				 i_9 => i_A(29),
				 i_10 => i_A(30),
				 i_11 => i_A(31),
				 i_12 => w_fill,
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(20));
	
	u_myMUX_bit19: myMUX32_1
	port map (i_0 => i_A(19),
				 i_1 => i_A(20),
				 i_2 => i_A(21),
				 i_3 => i_A(22),
				 i_4 => i_A(23),
				 i_5 => i_A(24),
				 i_6 => i_A(25),
				 i_7 => i_A(26),
				 i_8 => i_A(27),
				 i_9 => i_A(28),
				 i_10 => i_A(29),
				 i_11 => i_A(30),
				 i_12 => i_A(31),
				 i_13 => w_fill,
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(19));
	
	u_myMUX_bit18: myMUX32_1
	port map (i_0 => i_A(18),
				 i_1 => i_A(19),
				 i_2 => i_A(20),
				 i_3 => i_A(21),
				 i_4 => i_A(22),
				 i_5 => i_A(23),
				 i_6 => i_A(24),
				 i_7 => i_A(25),
				 i_8 => i_A(26),
				 i_9 => i_A(27),
				 i_10 => i_A(28),
				 i_11 => i_A(29),
				 i_12 => i_A(30),
				 i_13 => i_A(31),
				 i_14 => w_fill,
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(18));
	
	u_myMUX_bit17: myMUX32_1
	port map (i_0 => i_A(17),
				 i_1 => i_A(18),
				 i_2 => i_A(19),
				 i_3 => i_A(20),
				 i_4 => i_A(21),
				 i_5 => i_A(22),
				 i_6 => i_A(23),
				 i_7 => i_A(24),
				 i_8 => i_A(25),
				 i_9 => i_A(26),
				 i_10 => i_A(27),
				 i_11 => i_A(28),
				 i_12 => i_A(29),
				 i_13 => i_A(30),
				 i_14 => i_A(31),
				 i_15 => w_fill,
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(17));
	
	u_myMUX_bit16: myMUX32_1
	port map (i_0 => i_A(16),
				 i_1 => i_A(17),
				 i_2 => i_A(18),
				 i_3 => i_A(19),
				 i_4 => i_A(20),
				 i_5 => i_A(21),
				 i_6 => i_A(22),
				 i_7 => i_A(23),
				 i_8 => i_A(24),
				 i_9 => i_A(25),
				 i_10 => i_A(26),
				 i_11 => i_A(27),
				 i_12 => i_A(28),
				 i_13 => i_A(29),
				 i_14 => i_A(30),
				 i_15 => i_A(31),
				 i_16 => w_fill,
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(16));
				 
	u_myMUX_bit15: myMUX32_1
	port map (i_0 => i_A(15),
				 i_1 => i_A(16),
				 i_2 => i_A(17),
				 i_3 => i_A(18),
				 i_4 => i_A(19),
				 i_5 => i_A(20),
				 i_6 => i_A(21),
				 i_7 => i_A(22),
				 i_8 => i_A(23),
				 i_9 => i_A(24),
				 i_10 => i_A(25),
				 i_11 => i_A(26),
				 i_12 => i_A(27),
				 i_13 => i_A(28),
				 i_14 => i_A(29),
				 i_15 => i_A(30),
				 i_16 => i_A(31),
				 i_17 => w_fill,
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(15));
	
	u_myMUX_bit14: myMUX32_1
	port map (i_0 => i_A(14),
				 i_1 => i_A(15),
				 i_2 => i_A(16),
				 i_3 => i_A(17),
				 i_4 => i_A(18),
				 i_5 => i_A(19),
				 i_6 => i_A(20),
				 i_7 => i_A(21),
				 i_8 => i_A(22),
				 i_9 => i_A(23),
				 i_10 => i_A(24),
				 i_11 => i_A(25),
				 i_12 => i_A(26),
				 i_13 => i_A(27),
				 i_14 => i_A(28),
				 i_15 => i_A(29),
				 i_16 => i_A(30),
				 i_17 => i_A(31),
				 i_18 => w_fill,
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(14));
	
	u_myMUX_bit13: myMUX32_1
	port map (i_0 => i_A(13),
				 i_1 => i_A(14),
				 i_2 => i_A(15),
				 i_3 => i_A(16),
				 i_4 => i_A(17),
				 i_5 => i_A(18),
				 i_6 => i_A(19),
				 i_7 => i_A(20),
				 i_8 => i_A(21),
				 i_9 => i_A(22),
				 i_10 => i_A(23),
				 i_11 => i_A(24),
				 i_12 => i_A(25),
				 i_13 => i_A(26),
				 i_14 => i_A(27),
				 i_15 => i_A(28),
				 i_16 => i_A(29),
				 i_17 => i_A(30),
				 i_18 => i_A(31),
				 i_19 => w_fill,
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(13));
	
	u_myMUX_bit12: myMUX32_1
	port map (i_0 => i_A(12),
				 i_1 => i_A(13),
				 i_2 => i_A(14),
				 i_3 => i_A(15),
				 i_4 => i_A(16),
				 i_5 => i_A(17),
				 i_6 => i_A(18),
				 i_7 => i_A(19),
				 i_8 => i_A(20),
				 i_9 => i_A(21),
				 i_10 => i_A(22),
				 i_11 => i_A(23),
				 i_12 => i_A(24),
				 i_13 => i_A(25),
				 i_14 => i_A(26),
				 i_15 => i_A(27),
				 i_16 => i_A(28),
				 i_17 => i_A(29),
				 i_18 => i_A(30),
				 i_19 => i_A(31),
				 i_20 => w_fill,
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(12));
	
	u_myMUX_bit11: myMUX32_1
	port map (i_0 => i_A(11),
				 i_1 => i_A(12),
				 i_2 => i_A(13),
				 i_3 => i_A(14),
				 i_4 => i_A(15),
				 i_5 => i_A(16),
				 i_6 => i_A(17),
				 i_7 => i_A(18),
				 i_8 => i_A(19),
				 i_9 => i_A(20),
				 i_10 => i_A(21),
				 i_11 => i_A(22),
				 i_12 => i_A(23),
				 i_13 => i_A(24),
				 i_14 => i_A(25),
				 i_15 => i_A(26),
				 i_16 => i_A(27),
				 i_17 => i_A(28),
				 i_18 => i_A(29),
				 i_19 => i_A(30),
				 i_20 => i_A(31),
				 i_21 => w_fill,
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(11));
	
	u_myMUX_bit10: myMUX32_1
	port map (i_0 => i_A(10),
				 i_1 => i_A(11),
				 i_2 => i_A(12),
				 i_3 => i_A(13),
				 i_4 => i_A(14),
				 i_5 => i_A(15),
				 i_6 => i_A(16),
				 i_7 => i_A(17),
				 i_8 => i_A(18),
				 i_9 => i_A(19),
				 i_10 => i_A(20),
				 i_11 => i_A(21),
				 i_12 => i_A(22),
				 i_13 => i_A(23),
				 i_14 => i_A(24),
				 i_15 => i_A(25),
				 i_16 => i_A(26),
				 i_17 => i_A(27),
				 i_18 => i_A(28),
				 i_19 => i_A(29),
				 i_20 => i_A(30),
				 i_21 => i_A(31),
				 i_22 => w_fill,
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(10));
	
	u_myMUX_bit9: myMUX32_1
	port map (i_0 => i_A(9),
				 i_1 => i_A(10),
				 i_2 => i_A(11),
				 i_3 => i_A(12),
				 i_4 => i_A(13),
				 i_5 => i_A(14),
				 i_6 => i_A(15),
				 i_7 => i_A(16),
				 i_8 => i_A(17),
				 i_9 => i_A(18),
				 i_10 => i_A(19),
				 i_11 => i_A(20),
				 i_12 => i_A(21),
				 i_13 => i_A(22),
				 i_14 => i_A(23),
				 i_15 => i_A(24),
				 i_16 => i_A(25),
				 i_17 => i_A(26),
				 i_18 => i_A(27),
				 i_19 => i_A(28),
				 i_20 => i_A(29),
				 i_21 => i_A(30),
				 i_22 => i_A(31),
				 i_23 => w_fill,
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(9));
	
	u_myMUX_bit8: myMUX32_1
	port map (i_0 => i_A(8),
				 i_1 => i_A(9),
				 i_2 => i_A(10),
				 i_3 => i_A(11),
				 i_4 => i_A(12),
				 i_5 => i_A(13),
				 i_6 => i_A(14),
				 i_7 => i_A(15),
				 i_8 => i_A(16),
				 i_9 => i_A(17),
				 i_10 => i_A(18),
				 i_11 => i_A(19),
				 i_12 => i_A(20),
				 i_13 => i_A(21),
				 i_14 => i_A(22),
				 i_15 => i_A(23),
				 i_16 => i_A(24),
				 i_17 => i_A(25),
				 i_18 => i_A(26),
				 i_19 => i_A(27),
				 i_20 => i_A(28),
				 i_21 => i_A(29),
				 i_22 => i_A(30),
				 i_23 => i_A(31),
				 i_24 => w_fill,
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(8));
	
	u_myMUX_bit7: myMUX32_1
	port map (i_0 => i_A(7),
				 i_1 => i_A(8),
				 i_2 => i_A(9),
				 i_3 => i_A(10),
				 i_4 => i_A(11),
				 i_5 => i_A(12),
				 i_6 => i_A(13),
				 i_7 => i_A(14),
				 i_8 => i_A(15),
				 i_9 => i_A(16),
				 i_10 => i_A(17),
				 i_11 => i_A(18),
				 i_12 => i_A(19),
				 i_13 => i_A(20),
				 i_14 => i_A(21),
				 i_15 => i_A(22),
				 i_16 => i_A(23),
				 i_17 => i_A(24),
				 i_18 => i_A(25),
				 i_19 => i_A(26),
				 i_20 => i_A(27),
				 i_21 => i_A(28),
				 i_22 => i_A(29),
				 i_23 => i_A(30),
				 i_24 => i_A(31),
				 i_25 => w_fill,
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(7));
	
	u_myMUX_bit6: myMUX32_1
	port map (i_0 => i_A(6),
				 i_1 => i_A(7),
				 i_2 => i_A(8),
				 i_3 => i_A(9),
				 i_4 => i_A(10),
				 i_5 => i_A(11),
				 i_6 => i_A(12),
				 i_7 => i_A(13),
				 i_8 => i_A(14),
				 i_9 => i_A(15),
				 i_10 => i_A(16),
				 i_11 => i_A(17),
				 i_12 => i_A(18),
				 i_13 => i_A(19),
				 i_14 => i_A(20),
				 i_15 => i_A(21),
				 i_16 => i_A(22),
				 i_17 => i_A(23),
				 i_18 => i_A(24),
				 i_19 => i_A(25),
				 i_20 => i_A(26),
				 i_21 => i_A(27),
				 i_22 => i_A(28),
				 i_23 => i_A(29),
				 i_24 => i_A(30),
				 i_25 => i_A(31),
				 i_26 => w_fill,
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(6));
	
	u_myMUX_bit5: myMUX32_1
	port map (i_0 => i_A(5),
				 i_1 => i_A(6),
				 i_2 => i_A(7),
				 i_3 => i_A(8),
				 i_4 => i_A(9),
				 i_5 => i_A(10),
				 i_6 => i_A(11),
				 i_7 => i_A(12),
				 i_8 => i_A(13),
				 i_9 => i_A(14),
				 i_10 => i_A(15),
				 i_11 => i_A(16),
				 i_12 => i_A(17),
				 i_13 => i_A(18),
				 i_14 => i_A(19),
				 i_15 => i_A(20),
				 i_16 => i_A(21),
				 i_17 => i_A(22),
				 i_18 => i_A(23),
				 i_19 => i_A(24),
				 i_20 => i_A(25),
				 i_21 => i_A(26),
				 i_22 => i_A(27),
				 i_23 => i_A(28),
				 i_24 => i_A(29),
				 i_25 => i_A(30),
				 i_26 => i_A(31),
				 i_27 => w_fill,
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(5));
	
	u_myMUX_bit4: myMUX32_1
	port map (i_0 => i_A(4),
				 i_1 => i_A(5),
				 i_2 => i_A(6),
				 i_3 => i_A(7),
				 i_4 => i_A(8),
				 i_5 => i_A(9),
				 i_6 => i_A(10),
				 i_7 => i_A(11),
				 i_8 => i_A(12),
				 i_9 => i_A(13),
				 i_10 => i_A(14),
				 i_11 => i_A(15),
				 i_12 => i_A(16),
				 i_13 => i_A(17),
				 i_14 => i_A(18),
				 i_15 => i_A(19),
				 i_16 => i_A(20),
				 i_17 => i_A(21),
				 i_18 => i_A(22),
				 i_19 => i_A(23),
				 i_20 => i_A(24),
				 i_21 => i_A(25),
				 i_22 => i_A(26),
				 i_23 => i_A(27),
				 i_24 => i_A(28),
				 i_25 => i_A(29),
				 i_26 => i_A(30),
				 i_27 => i_A(31),
				 i_28 => w_fill,
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(4));
	
	u_myMUX_bit3: myMUX32_1
	port map (i_0 => i_A(3),
				 i_1 => i_A(4),
				 i_2 => i_A(5),
				 i_3 => i_A(6),
				 i_4 => i_A(7),
				 i_5 => i_A(8),
				 i_6 => i_A(9),
				 i_7 => i_A(10),
				 i_8 => i_A(11),
				 i_9 => i_A(12),
				 i_10 => i_A(13),
				 i_11 => i_A(14),
				 i_12 => i_A(15),
				 i_13 => i_A(16),
				 i_14 => i_A(17),
				 i_15 => i_A(18),
				 i_16 => i_A(19),
				 i_17 => i_A(20),
				 i_18 => i_A(21),
				 i_19 => i_A(22),
				 i_20 => i_A(23),
				 i_21 => i_A(24),
				 i_22 => i_A(25),
				 i_23 => i_A(26),
				 i_24 => i_A(27),
				 i_25 => i_A(28),
				 i_26 => i_A(29),
				 i_27 => i_A(30),
				 i_28 => i_A(31),
				 i_29 => w_fill,
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(3));
	
	u_myMUX_bit2: myMUX32_1
	port map (i_0 => i_A(2),
				 i_1 => i_A(3),
				 i_2 => i_A(4),
				 i_3 => i_A(5),
				 i_4 => i_A(6),
				 i_5 => i_A(7),
				 i_6 => i_A(8),
				 i_7 => i_A(9),
				 i_8 => i_A(10),
				 i_9 => i_A(11),
				 i_10 => i_A(12),
				 i_11 => i_A(13),
				 i_12 => i_A(14),
				 i_13 => i_A(15),
				 i_14 => i_A(16),
				 i_15 => i_A(17),
				 i_16 => i_A(18),
				 i_17 => i_A(19),
				 i_18 => i_A(20),
				 i_19 => i_A(21),
				 i_20 => i_A(22),
				 i_21 => i_A(23),
				 i_22 => i_A(24),
				 i_23 => i_A(25),
				 i_24 => i_A(26),
				 i_25 => i_A(27),
				 i_26 => i_A(28),
				 i_27 => i_A(29),
				 i_28 => i_A(30),
				 i_29 => i_A(31),
				 i_30 => w_fill,
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(2));
	
	u_myMUX_bit1: myMUX32_1
	port map (i_0 => i_A(1),
				 i_1 => i_A(2),
				 i_2 => i_A(3),
				 i_3 => i_A(4),
				 i_4 => i_A(5),
				 i_5 => i_A(6),
				 i_6 => i_A(7),
				 i_7 => i_A(8),
				 i_8 => i_A(9),
				 i_9 => i_A(10),
				 i_10 => i_A(11),
				 i_11 => i_A(12),
				 i_12 => i_A(13),
				 i_13 => i_A(14),
				 i_14 => i_A(15),
				 i_15 => i_A(16),
				 i_16 => i_A(17),
				 i_17 => i_A(18),
				 i_18 => i_A(19),
				 i_19 => i_A(20),
				 i_20 => i_A(21),
				 i_21 => i_A(22),
				 i_22 => i_A(23),
				 i_23 => i_A(24),
				 i_24 => i_A(25),
				 i_25 => i_A(26),
				 i_26 => i_A(27),
				 i_27 => i_A(28),
				 i_28 => i_A(29),
				 i_29 => i_A(30),
				 i_30 => i_A(31),
				 i_31 => w_fill,
				 i_S => i_SA,
				 o_Z => o_Z(1));
				 
	u_myMUX_bit0: myMUX32_1
	port map (i_0 => i_A(0),
				 i_1 => i_A(1),
				 i_2 => i_A(2),
				 i_3 => i_A(3),
				 i_4 => i_A(4),
				 i_5 => i_A(5),
				 i_6 => i_A(6),
				 i_7 => i_A(7),
				 i_8 => i_A(8),
				 i_9 => i_A(9),
				 i_10 => i_A(10),
				 i_11 => i_A(11),
				 i_12 => i_A(12),
				 i_13 => i_A(13),
				 i_14 => i_A(14),
				 i_15 => i_A(15),
				 i_16 => i_A(16),
				 i_17 => i_A(17),
				 i_18 => i_A(18),
				 i_19 => i_A(19),
				 i_20 => i_A(20),
				 i_21 => i_A(21),
				 i_22 => i_A(22),
				 i_23 => i_A(23),
				 i_24 => i_A(24),
				 i_25 => i_A(25),
				 i_26 => i_A(26),
				 i_27 => i_A(27),
				 i_28 => i_A(28),
				 i_29 => i_A(29),
				 i_30 => i_A(30),
				 i_31 => i_A(31),
				 i_S => i_SA,
				 o_Z => o_Z(0));
end a_RIGHT_SHIFT;