--| Test32_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:10:14
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test32_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test32_Reg_COMBINED;

architecture a_Test32_Reg_COMBINED of Test32_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 466) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 466) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100");--  465 - 1860

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000011000010011011111", --    2 -    8
      "00101000000000100001010111011001", --    3 -   12
      "00101100000000110000100011111011", --    4 -   16
      "00000000010000000010000000000100", --    5 -   20
      "00000000010000000010100000100011", --    6 -   24
      "00000000010001010011000000100000", --    7 -   28
      "00000000100001000011100000101010", --    8 -   32
      "00000000111001000100000000100001", --    9 -   36
      "00101100000010011011110101111111", --   10 -   40
      "00000001000000000101000000100111", --   11 -   44
      "00000001010010010101100000100100", --   12 -   48
      "00100100111011000110110011101000", --   13 -   52
      "00100000101011010111110111100101", --   14 -   56
      "00101000110011100001000110000100", --   15 -   60
      "00110100101011110101010110011111", --   16 -   64
      "00000001000010001000000000100101", --   17 -   68
      "00000001000000001000100000100010", --   18 -   72
      "00000001111011011001000000100001", --   19 -   76
      "00000000111000011001100000000100", --   20 -   80
      "00000000101011101010000000100000", --   21 -   84
      "00000010000100111010100000100000", --   22 -   88
      "00000000000000000000000000000000", --   23 -   92
      "00100000100101101000110010110101", --   24 -   96
      "00000000000000000000000000000000", --   25 -  100
      "00000010010010111011100000100010", --   26 -  104
      "00000001100000001100000000100110", --   27 -  108
      "00100110100110010110000001100110", --   28 -  112
      "10101100000100010000001100101100", --   29 -  116
      "00110010100110101011001011011010", --   30 -  120
      "00000000000000000000000000000000", --   31 -  124
      "10101100000110000000001100110000", --   32 -  128
      "10101100000101110000001100110100", --   33 -  132
      "00100110110110111010000010110001", --   34 -  136
      "10101100000110100000001100111000", --   35 -  140
      "00000000000000000000000000000000", --   36 -  144
      "00000011011010001110000000000110", --   37 -  148
      "00111100000111011101000111110000", --   38 -  152
      "10101100000111000000001100111100", --   39 -  156
      "00101000011111101011011110100110", --   40 -  160
      "00101010110000101010010111101111", --   41 -  164
      "10101100000000100000001101000000", --   42 -  168
      "00111100000010100111001101000100", --   43 -  172
      "00000011000111010100100000100011", --   44 -  176
      "00000000000000000000000000000000", --   45 -  180
      "00000011001011000011000000000110", --   46 -  184
      "10101100000010000000001101000100", --   47 -  188
      "00000000110101010111100000100111", --   48 -  192
      "10101100000101010000001101001000", --   49 -  196
      "10101100000011110000001101001100", --   50 -  200
      "00000001010011010000100000101010", --   51 -  204
      "00000001001111100100100000100001", --   52 -  208
      "10101100000010000000001101010000", --   53 -  212
      "00000000000000000000000000000000", --   54 -  216
      "00000000000000000000000000000000", --   55 -  220
      "00000000000000010011100011000000", --   56 -  224
      "00000000000000010010101001000011", --   57 -  228
      "00100001001011101100101101101010", --   58 -  232
      "10101100000001110000001101010100", --   59 -  236
      "10101100000001010000001101011000", --   60 -  240
      "10101100000011100000001101011100", --   61 -  244
      "10101100000010010000001101100000", --   62 -  248
      "00100011111111111111111111111111", --   63 -  252
      "00011111111000001111111111000010", --   64 -  256
      "00010000000000000000000110010000", --   65 -  260
      "00111100000111100000001111100111", --   66 -  264
      "00111100000111110000001111100111", --   67 -  268
      "00000000000111101111010000000010", --   68 -  272
      "00000000000111111111110000000010", --   69 -  276
      "00111100000000011000010011011111", --   70 -  280
      "00111100000011111000010011011111", --   71 -  284
      "00101000000000100001010111011001", --   72 -  288
      "00101000000100000001010111011001", --   73 -  292
      "00101100000000110000100011111011", --   74 -  296
      "00101100000100010000100011111011", --   75 -  300
      "00000000010000000010000000000100", --   76 -  304
      "00000010000000001001000000000100", --   77 -  308
      "00000000010000000010100000100011", --   78 -  312
      "00000010000000001001100000100011", --   79 -  316
      "00000000010001010011000000100000", --   80 -  320
      "00000010000100111010000000100000", --   81 -  324
      "00000000100001000011100000101010", --   82 -  328
      "00000010010100101010100000101010", --   83 -  332
      "00000000111001000100000000100001", --   84 -  336
      "00000010101100101011000000100001", --   85 -  340
      "00101100000010011011110101111111", --   86 -  344
      "00101100000101111011110101111111", --   87 -  348
      "00000001000000000101000000100111", --   88 -  352
      "00000010110000001100000000100111", --   89 -  356
      "00000001010010010101100000100100", --   90 -  360
      "00000011000101111100100000100100", --   91 -  364
      "00100100111011000110110011101000", --   92 -  368
      "00100110101110100110110011101000", --   93 -  372
      "00100000101011010111110111100101", --   94 -  376
      "00100010011110110111110111100101", --   95 -  380
      "00101000110011100001000110000100", --   96 -  384
      "00101010100111000001000110000100", --   97 -  388
      "00110100101000100101010110011111", --   98 -  392
      "00110110011100000101010110011111", --   99 -  396
      "00000001000010000101000000100101", --  100 -  400
      "00000010110101101100000000100101", --  101 -  404
      "00000001000000000100100000100010", --  102 -  408
      "00000010110000001011100000100010", --  103 -  412
      "00000000010011010011000000100001", --  104 -  416
      "00000010000110111010000000100001", --  105 -  420
      "00000000111000010001000000000100", --  106 -  424
      "00000010101011111000000000000100", --  107 -  428
      "00000000101011100000100000100000", --  108 -  432
      "00000010011111000111100000100000", --  109 -  436
      "00000001010000100011100000100000", --  110 -  440
      "00000011000100001010100000100000", --  111 -  444
      "00000000000000000000000000000000", --  112 -  448
      "00000000000000000000000000000000", --  113 -  452
      "00100000100001011000110010110101", --  114 -  456
      "00100010010100111000110010110101", --  115 -  460
      "00000000000000000000000000000000", --  116 -  464
      "00000000000000000000000000000000", --  117 -  468
      "00000000110010110111000000100010", --  118 -  472
      "00000010100110011110000000100010", --  119 -  476
      "00000001100000000101000000100110", --  120 -  480
      "00000011010000001100000000100110", --  121 -  484
      "00100100001000100110000001100110", --  122 -  488
      "00100101111100000110000001100110", --  123 -  492
      "00010101001101110000000011001000", --  124 -  496
      "10101100000010010000001100101100", --  125 -  500
      "00110000001001001011001011011010", --  126 -  504
      "00110001111100101011001011011010", --  127 -  508
      "00000000000000000000000000000000", --  128 -  512
      "00000000000000000000000000000000", --  129 -  516
      "00010101010110000000000011000010", --  130 -  520
      "10101100000010100000001100110000", --  131 -  524
      "00010101110111000000000011000000", --  132 -  528
      "10101100000011100000001100110100", --  133 -  532
      "00100100101001101010000010110001", --  134 -  536
      "00100110011101001010000010110001", --  135 -  540
      "00010100100100100000000010111100", --  136 -  544
      "10101100000001000000001100111000", --  137 -  548
      "00000000000000000000000000000000", --  138 -  552
      "00000000000000000000000000000000", --  139 -  556
      "00000000110010000101100000000110", --  140 -  560
      "00000010100101101100100000000110", --  141 -  564
      "00111100000010011101000111110000", --  142 -  568
      "00111100000101111101000111110000", --  143 -  572
      "00010101011110010000000010110100", --  144 -  576
      "10101100000010110000001100111100", --  145 -  580
      "00101000011000011011011110100110", --  146 -  584
      "00101010001011111011011110100110", --  147 -  588
      "00101000101011101010010111101111", --  148 -  592
      "00101010011111001010010111101111", --  149 -  596
      "00010101110111000000000010101110", --  150 -  600
      "10101100000011100000001101000000", --  151 -  604
      "00111100000001000111001101000100", --  152 -  608
      "00111100000100100111001101000100", --  153 -  612
      "00000001010010010011000000100011", --  154 -  616
      "00000011000101111010000000100011", --  155 -  620
      "00000000000000000000000000000000", --  156 -  624
      "00000000000000000000000000000000", --  157 -  628
      "00000000010011000101100000000110", --  158 -  632
      "00000010000110101100100000000110", --  159 -  636
      "00010101000101100000000010100100", --  160 -  640
      "10101100000010000000001101000100", --  161 -  644
      "00000001011001110001100000100111", --  162 -  648
      "00000011001101011000100000100111", --  163 -  652
      "00010100111101010000000010100000", --  164 -  656
      "10101100000001110000001101001000", --  165 -  660
      "00010100011100010000000010011110", --  166 -  664
      "10101100000000110000001101001100", --  167 -  668
      "00000000100011010010100000101010", --  168 -  672
      "00000010010110111001100000101010", --  169 -  676
      "00000000110000010011000000100001", --  170 -  680
      "00000010100011111010000000100001", --  171 -  684
      "00010101000101100000000010011000", --  172 -  688
      "10101100000010000000001101010000", --  173 -  692
      "00000000000000000000000000000000", --  174 -  696
      "00000000000000000000000000000000", --  175 -  700
      "00000000000000000000000000000000", --  176 -  704
      "00000000000000000000000000000000", --  177 -  708
      "00000000000001010111000011000000", --  178 -  712
      "00000000000100111110000011000000", --  179 -  716
      "00000000000001010101001001000011", --  180 -  720
      "00000000000100111100001001000011", --  181 -  724
      "00100000110010011100101101101010", --  182 -  728
      "00100010100101111100101101101010", --  183 -  732
      "00010101110111000000000010001100", --  184 -  736
      "10101100000011100000001101010100", --  185 -  740
      "00010101010110000000000010001010", --  186 -  744
      "10101100000010100000001101011000", --  187 -  748
      "00010101001101110000000010001000", --  188 -  752
      "10101100000010010000001101011100", --  189 -  756
      "00010100110101000000000010000110", --  190 -  760
      "10101100000001100000001101100000", --  191 -  764
      "00100011110111011111111100000110", --  192 -  768
      "00010011101000000000000000011000", --  193 -  772
      "00100011110111011111111000001100", --  194 -  776
      "00010011101000000000000000010110", --  195 -  780
      "00100011110111011111110100010010", --  196 -  784
      "00010011101000000000000000010100", --  197 -  788
      "00100011110111101111111111111111", --  198 -  792
      "00100011111111111111111111111111", --  199 -  796
      "00010111110111110000000001111100", --  200 -  800
      "00011111111000001111111101111101", --  201 -  804
      "00010000000000000000000100000111", --  202 -  808
      "00000000000000000000000000000000", --  203 -  812
      "00000000000000000000000000000000", --  204 -  816
      "00000000000000000000000000000000", --  205 -  820
      "00000000000000000000000000000000", --  206 -  824
      "00000000000000000000000000000000", --  207 -  828
      "00000000000000000000000000000000", --  208 -  832
      "00000000000000000000000000000000", --  209 -  836
      "00000000000000000000000000000000", --  210 -  840
      "00000000000000000000000000000000", --  211 -  844
      "00000000000000000000000000000000", --  212 -  848
      "00000000000000000000000000000000", --  213 -  852
      "00000000000000000000000000000000", --  214 -  856
      "00000000000000000000000000000000", --  215 -  860
      "00000000000000000000000000000000", --  216 -  864
      "10001100000111010000011010111000", --  217 -  868
      "00011111101000000000000000000011", --  218 -  872
      "00100000000111010000000000111100", --  219 -  876
      "00010000000000000000000000000010", --  220 -  880
      "00100000000111010000000000000000", --  221 -  884
      "00010100001011110000000001100110", --  222 -  888
      "10101111101000010000011001000000", --  223 -  892
      "10001100000111010000011010111000", --  224 -  896
      "00011111101000000000000000000011", --  225 -  900
      "00100000000111010000000000111100", --  226 -  904
      "00010000000000000000000000000010", --  227 -  908
      "00100000000111010000000000000000", --  228 -  912
      "00010100010100000000000001011111", --  229 -  916
      "10101111101000100000011001000100", --  230 -  920
      "10001100000111010000011010111000", --  231 -  924
      "00011111101000000000000000000011", --  232 -  928
      "00100000000111010000000000111100", --  233 -  932
      "00010000000000000000000000000010", --  234 -  936
      "00100000000111010000000000000000", --  235 -  940
      "00010100011100010000000001011000", --  236 -  944
      "10101111101000110000011001001000", --  237 -  948
      "10001100000111010000011010111000", --  238 -  952
      "00011111101000000000000000000011", --  239 -  956
      "00100000000111010000000000111100", --  240 -  960
      "00010000000000000000000000000010", --  241 -  964
      "00100000000111010000000000000000", --  242 -  968
      "00010100100100100000000001010001", --  243 -  972
      "10101111101001000000011001001100", --  244 -  976
      "10001100000111010000011010111000", --  245 -  980
      "00011111101000000000000000000011", --  246 -  984
      "00100000000111010000000000111100", --  247 -  988
      "00010000000000000000000000000010", --  248 -  992
      "00100000000111010000000000000000", --  249 -  996
      "00010100101100110000000001001010", --  250 - 1000
      "10101111101001010000011001010000", --  251 - 1004
      "10001100000111010000011010111000", --  252 - 1008
      "00011111101000000000000000000011", --  253 - 1012
      "00100000000111010000000000111100", --  254 - 1016
      "00010000000000000000000000000010", --  255 - 1020
      "00100000000111010000000000000000", --  256 - 1024
      "00010100110101000000000001000011", --  257 - 1028
      "10101111101001100000011001010100", --  258 - 1032
      "10001100000111010000011010111000", --  259 - 1036
      "00011111101000000000000000000011", --  260 - 1040
      "00100000000111010000000000111100", --  261 - 1044
      "00010000000000000000000000000010", --  262 - 1048
      "00100000000111010000000000000000", --  263 - 1052
      "00010100111101010000000000111100", --  264 - 1056
      "10101111101001110000011001011000", --  265 - 1060
      "10001100000111010000011010111000", --  266 - 1064
      "00011111101000000000000000000011", --  267 - 1068
      "00100000000111010000000000111100", --  268 - 1072
      "00010000000000000000000000000010", --  269 - 1076
      "00100000000111010000000000000000", --  270 - 1080
      "00010101000101100000000000110101", --  271 - 1084
      "10101111101010000000011001011100", --  272 - 1088
      "10001100000111010000011010111000", --  273 - 1092
      "00011111101000000000000000000011", --  274 - 1096
      "00100000000111010000000000111100", --  275 - 1100
      "00010000000000000000000000000010", --  276 - 1104
      "00100000000111010000000000000000", --  277 - 1108
      "00010101001101110000000000101110", --  278 - 1112
      "10101111101010010000011001100000", --  279 - 1116
      "10001100000111010000011010111000", --  280 - 1120
      "00011111101000000000000000000011", --  281 - 1124
      "00100000000111010000000000111100", --  282 - 1128
      "00010000000000000000000000000010", --  283 - 1132
      "00100000000111010000000000000000", --  284 - 1136
      "00010101010110000000000000100111", --  285 - 1140
      "10101111101010100000011001100100", --  286 - 1144
      "10001100000111010000011010111000", --  287 - 1148
      "00011111101000000000000000000011", --  288 - 1152
      "00100000000111010000000000111100", --  289 - 1156
      "00010000000000000000000000000010", --  290 - 1160
      "00100000000111010000000000000000", --  291 - 1164
      "00010101011110010000000000100000", --  292 - 1168
      "10101111101010110000011001101000", --  293 - 1172
      "10001100000111010000011010111000", --  294 - 1176
      "00011111101000000000000000000011", --  295 - 1180
      "00100000000111010000000000111100", --  296 - 1184
      "00010000000000000000000000000010", --  297 - 1188
      "00100000000111010000000000000000", --  298 - 1192
      "00010101100110100000000000011001", --  299 - 1196
      "10101111101011000000011001101100", --  300 - 1200
      "10001100000111010000011010111000", --  301 - 1204
      "00011111101000000000000000000011", --  302 - 1208
      "00100000000111010000000000111100", --  303 - 1212
      "00010000000000000000000000000010", --  304 - 1216
      "00100000000111010000000000000000", --  305 - 1220
      "00010101101110110000000000010010", --  306 - 1224
      "10101111101011010000011001110000", --  307 - 1228
      "10001100000111010000011010111000", --  308 - 1232
      "00011111101000000000000000000011", --  309 - 1236
      "00100000000111010000000000111100", --  310 - 1240
      "00010000000000000000000000000010", --  311 - 1244
      "00100000000111010000000000000000", --  312 - 1248
      "00010101110111000000000000001011", --  313 - 1252
      "10101111101011100000011001110100", --  314 - 1256
      "10001100000111010000011010111000", --  315 - 1260
      "00011111101000000000000000000011", --  316 - 1264
      "00100000000111010000000000111100", --  317 - 1268
      "00010000000000000000000000000010", --  318 - 1272
      "00100000000111010000000000000000", --  319 - 1276
      "00010111110111110000000000000100", --  320 - 1280
      "10101111101111100000011001111000", --  321 - 1284
      "10101100000111010000011010111000", --  322 - 1288
      "00010000000000001111111110000011", --  323 - 1292
      "10001100000111010000011010111000", --  324 - 1296
      "10001111101000010000011001000000", --  325 - 1300
      "10001100000111010000011010111000", --  326 - 1304
      "10001111101011110000011001000000", --  327 - 1308
      "00010100001011111111111111111100", --  328 - 1312
      "10001100000111010000011010111000", --  329 - 1316
      "10001111101000100000011001000100", --  330 - 1320
      "10001100000111010000011010111000", --  331 - 1324
      "10001111101100000000011001000100", --  332 - 1328
      "00010100010100001111111111111100", --  333 - 1332
      "10001100000111010000011010111000", --  334 - 1336
      "10001111101000110000011001001000", --  335 - 1340
      "10001100000111010000011010111000", --  336 - 1344
      "10001111101100010000011001001000", --  337 - 1348
      "00010100011100011111111111111100", --  338 - 1352
      "10001100000111010000011010111000", --  339 - 1356
      "10001111101001000000011001001100", --  340 - 1360
      "10001100000111010000011010111000", --  341 - 1364
      "10001111101100100000011001001100", --  342 - 1368
      "00010100100100101111111111111100", --  343 - 1372
      "10001100000111010000011010111000", --  344 - 1376
      "10001111101001010000011001010000", --  345 - 1380
      "10001100000111010000011010111000", --  346 - 1384
      "10001111101100110000011001010000", --  347 - 1388
      "00010100101100111111111111111100", --  348 - 1392
      "10001100000111010000011010111000", --  349 - 1396
      "10001111101001100000011001010100", --  350 - 1400
      "10001100000111010000011010111000", --  351 - 1404
      "10001111101101000000011001010100", --  352 - 1408
      "00010100110101001111111111111100", --  353 - 1412
      "10001100000111010000011010111000", --  354 - 1416
      "10001111101001110000011001011000", --  355 - 1420
      "10001100000111010000011010111000", --  356 - 1424
      "10001111101101010000011001011000", --  357 - 1428
      "00010100111101011111111111111100", --  358 - 1432
      "10001100000111010000011010111000", --  359 - 1436
      "10001111101010000000011001011100", --  360 - 1440
      "10001100000111010000011010111000", --  361 - 1444
      "10001111101101100000011001011100", --  362 - 1448
      "00010101000101101111111111111100", --  363 - 1452
      "10001100000111010000011010111000", --  364 - 1456
      "10001111101010010000011001100000", --  365 - 1460
      "10001100000111010000011010111000", --  366 - 1464
      "10001111101101110000011001100000", --  367 - 1468
      "00010101001101111111111111111100", --  368 - 1472
      "10001100000111010000011010111000", --  369 - 1476
      "10001111101010100000011001100100", --  370 - 1480
      "10001100000111010000011010111000", --  371 - 1484
      "10001111101110000000011001100100", --  372 - 1488
      "00010101010110001111111111111100", --  373 - 1492
      "10001100000111010000011010111000", --  374 - 1496
      "10001111101010110000011001101000", --  375 - 1500
      "10001100000111010000011010111000", --  376 - 1504
      "10001111101110010000011001101000", --  377 - 1508
      "00010101011110011111111111111100", --  378 - 1512
      "10001100000111010000011010111000", --  379 - 1516
      "10001111101011000000011001101100", --  380 - 1520
      "10001100000111010000011010111000", --  381 - 1524
      "10001111101110100000011001101100", --  382 - 1528
      "00010101100110101111111111111100", --  383 - 1532
      "10001100000111010000011010111000", --  384 - 1536
      "10001111101011010000011001110000", --  385 - 1540
      "10001100000111010000011010111000", --  386 - 1544
      "10001111101110110000011001110000", --  387 - 1548
      "00010101101110111111111111111100", --  388 - 1552
      "10001100000111010000011010111000", --  389 - 1556
      "10001111101011100000011001110100", --  390 - 1560
      "10001100000111010000011010111000", --  391 - 1564
      "10001111101111000000011001110100", --  392 - 1568
      "00010101110111001111111111111100", --  393 - 1572
      "10001100000111010000011010111000", --  394 - 1576
      "10001111101111100000011001111000", --  395 - 1580
      "10001100000111010000011010111000", --  396 - 1584
      "10001111101111110000011001111000", --  397 - 1588
      "00010111110111111111111111111100", --  398 - 1592
      "00010000000000001111111100110111", --  399 - 1596
      "00000000000000000000000000000000", --  400 - 1600
      "00000000000000000000000000000000", --  401 - 1604
      "00000000000000000000000000000000", --  402 - 1608
      "00000000000000000000000000000000", --  403 - 1612
      "00000000000000000000000000000000", --  404 - 1616
      "00000000000000000000000000000000", --  405 - 1620
      "00000000000000000000000000000000", --  406 - 1624
      "00000000000000000000000000000000", --  407 - 1628
      "00000000000000000000000000000000", --  408 - 1632
      "00000000000000000000000000000000", --  409 - 1636
      "00000000000000000000000000000000", --  410 - 1640
      "00000000000000000000000000000000", --  411 - 1644
      "00000000000000000000000000000000", --  412 - 1648
      "00000000000000000000000000000000", --  413 - 1652
      "00000000000000000000000000000000", --  414 - 1656
      "00000000000000000000000000000000", --  415 - 1660
      "00000000000000000000000000000000", --  416 - 1664
      "00000000000000000000000000000000", --  417 - 1668
      "00000000000000000000000000000000", --  418 - 1672
      "00000000000000000000000000000000", --  419 - 1676
      "00000000000000000000000000000000", --  420 - 1680
      "00000000000000000000000000000000", --  421 - 1684
      "00000000000000000000000000000000", --  422 - 1688
      "00000000000000000000000000000000", --  423 - 1692
      "00000000000000000000000000000000", --  424 - 1696
      "00000000000000000000000000000000", --  425 - 1700
      "00000000000000000000000000000000", --  426 - 1704
      "00000000000000000000000000000000", --  427 - 1708
      "00000000000000000000000000000000", --  428 - 1712
      "00000000000000000000000000000000", --  429 - 1716
      "00000000000000000000001111100111", --  430 - 1720
      "00000000000000000000000000000000", --  431 - 1724
      "00000000000000000000000000000000", --  432 - 1728
      "00000000000000000000000000000000", --  433 - 1732
      "00000000000000000000000000000000", --  434 - 1736
      "00000000000000000000000000000000", --  435 - 1740
      "00000000000000000000000000000000", --  436 - 1744
      "00000000000000000000000000000000", --  437 - 1748
      "00000000000000000000000000000000", --  438 - 1752
      "00000000000000000000000000000000", --  439 - 1756
      "00000000000000000000000000000000", --  440 - 1760
      "00000000000000000000000000000000", --  441 - 1764
      "00000000000000000000000000000000", --  442 - 1768
      "00000000000000000000000000000000", --  443 - 1772
      "00000000000000000000000000000000", --  444 - 1776
      "00000000000000000000000000000000", --  445 - 1780
      "00000000000000000000000000000000", --  446 - 1784
      "00000000000000000000000000000000", --  447 - 1788
      "00000000000000000000000000000000", --  448 - 1792
      "00000000000000000000000000000000", --  449 - 1796
      "00000000000000000000000000000000", --  450 - 1800
      "00000000000000000000000000000000", --  451 - 1804
      "00000000000000000000000000000000", --  452 - 1808
      "00000000000000000000000000000000", --  453 - 1812
      "00000000000000000000000000000000", --  454 - 1816
      "00000000000000000000000000000000", --  455 - 1820
      "00000000000000000000000000000000", --  456 - 1824
      "00000000000000000000000000000000", --  457 - 1828
      "00000000000000000000000000000000", --  458 - 1832
      "00000000000000000000000000000000", --  459 - 1836
      "00000000000000000000000000000000", --  460 - 1840
      "00000000000000000000000000000000", --  461 - 1844
      "00000000000000000000000000000000", --  462 - 1848
      "00000000000000000000000000000000", --  463 - 1852
      "00000000000000000000000000000000", --  464 - 1856
      "00000000000000000000000000000000");--  465 - 1860

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000011000010011011111";
         f_reg(4) <= "00101000000000100001010111011001";
         f_reg(5) <= "00101100000000110000100011111011";
         f_reg(6) <= "00000000010000000010000000000100";
         f_reg(7) <= "00000000010000000010100000100011";
         f_reg(8) <= "00000000010001010011000000100000";
         f_reg(9) <= "00000000100001000011100000101010";
         f_reg(10) <= "00000000111001000100000000100001";
         f_reg(11) <= "00101100000010011011110101111111";
         f_reg(12) <= "00000001000000000101000000100111";
         f_reg(13) <= "00000001010010010101100000100100";
         f_reg(14) <= "00100100111011000110110011101000";
         f_reg(15) <= "00100000101011010111110111100101";
         f_reg(16) <= "00101000110011100001000110000100";
         f_reg(17) <= "00110100101011110101010110011111";
         f_reg(18) <= "00000001000010001000000000100101";
         f_reg(19) <= "00000001000000001000100000100010";
         f_reg(20) <= "00000001111011011001000000100001";
         f_reg(21) <= "00000000111000011001100000000100";
         f_reg(22) <= "00000000101011101010000000100000";
         f_reg(23) <= "00000010000100111010100000100000";
         f_reg(24) <= "00000000000000000000000000000000";
         f_reg(25) <= "00100000100101101000110010110101";
         f_reg(26) <= "00000000000000000000000000000000";
         f_reg(27) <= "00000010010010111011100000100010";
         f_reg(28) <= "00000001100000001100000000100110";
         f_reg(29) <= "00100110100110010110000001100110";
         f_reg(30) <= "10101100000100010000001100101100";
         f_reg(31) <= "00110010100110101011001011011010";
         f_reg(32) <= "00000000000000000000000000000000";
         f_reg(33) <= "10101100000110000000001100110000";
         f_reg(34) <= "10101100000101110000001100110100";
         f_reg(35) <= "00100110110110111010000010110001";
         f_reg(36) <= "10101100000110100000001100111000";
         f_reg(37) <= "00000000000000000000000000000000";
         f_reg(38) <= "00000011011010001110000000000110";
         f_reg(39) <= "00111100000111011101000111110000";
         f_reg(40) <= "10101100000111000000001100111100";
         f_reg(41) <= "00101000011111101011011110100110";
         f_reg(42) <= "00101010110000101010010111101111";
         f_reg(43) <= "10101100000000100000001101000000";
         f_reg(44) <= "00111100000010100111001101000100";
         f_reg(45) <= "00000011000111010100100000100011";
         f_reg(46) <= "00000000000000000000000000000000";
         f_reg(47) <= "00000011001011000011000000000110";
         f_reg(48) <= "10101100000010000000001101000100";
         f_reg(49) <= "00000000110101010111100000100111";
         f_reg(50) <= "10101100000101010000001101001000";
         f_reg(51) <= "10101100000011110000001101001100";
         f_reg(52) <= "00000001010011010000100000101010";
         f_reg(53) <= "00000001001111100100100000100001";
         f_reg(54) <= "10101100000010000000001101010000";
         f_reg(55) <= "00000000000000000000000000000000";
         f_reg(56) <= "00000000000000000000000000000000";
         f_reg(57) <= "00000000000000010011100011000000";
         f_reg(58) <= "00000000000000010010101001000011";
         f_reg(59) <= "00100001001011101100101101101010";
         f_reg(60) <= "10101100000001110000001101010100";
         f_reg(61) <= "10101100000001010000001101011000";
         f_reg(62) <= "10101100000011100000001101011100";
         f_reg(63) <= "10101100000010010000001101100000";
         f_reg(64) <= "00100011111111111111111111111111";
         f_reg(65) <= "00011111111000001111111111000010";
         f_reg(66) <= "00010000000000000000000110010000";
         f_reg(67) <= "00111100000111100000001111100111";
         f_reg(68) <= "00111100000111110000001111100111";
         f_reg(69) <= "00000000000111101111010000000010";
         f_reg(70) <= "00000000000111111111110000000010";
         f_reg(71) <= "00111100000000011000010011011111";
         f_reg(72) <= "00111100000011111000010011011111";
         f_reg(73) <= "00101000000000100001010111011001";
         f_reg(74) <= "00101000000100000001010111011001";
         f_reg(75) <= "00101100000000110000100011111011";
         f_reg(76) <= "00101100000100010000100011111011";
         f_reg(77) <= "00000000010000000010000000000100";
         f_reg(78) <= "00000010000000001001000000000100";
         f_reg(79) <= "00000000010000000010100000100011";
         f_reg(80) <= "00000010000000001001100000100011";
         f_reg(81) <= "00000000010001010011000000100000";
         f_reg(82) <= "00000010000100111010000000100000";
         f_reg(83) <= "00000000100001000011100000101010";
         f_reg(84) <= "00000010010100101010100000101010";
         f_reg(85) <= "00000000111001000100000000100001";
         f_reg(86) <= "00000010101100101011000000100001";
         f_reg(87) <= "00101100000010011011110101111111";
         f_reg(88) <= "00101100000101111011110101111111";
         f_reg(89) <= "00000001000000000101000000100111";
         f_reg(90) <= "00000010110000001100000000100111";
         f_reg(91) <= "00000001010010010101100000100100";
         f_reg(92) <= "00000011000101111100100000100100";
         f_reg(93) <= "00100100111011000110110011101000";
         f_reg(94) <= "00100110101110100110110011101000";
         f_reg(95) <= "00100000101011010111110111100101";
         f_reg(96) <= "00100010011110110111110111100101";
         f_reg(97) <= "00101000110011100001000110000100";
         f_reg(98) <= "00101010100111000001000110000100";
         f_reg(99) <= "00110100101000100101010110011111";
         f_reg(100) <= "00110110011100000101010110011111";
         f_reg(101) <= "00000001000010000101000000100101";
         f_reg(102) <= "00000010110101101100000000100101";
         f_reg(103) <= "00000001000000000100100000100010";
         f_reg(104) <= "00000010110000001011100000100010";
         f_reg(105) <= "00000000010011010011000000100001";
         f_reg(106) <= "00000010000110111010000000100001";
         f_reg(107) <= "00000000111000010001000000000100";
         f_reg(108) <= "00000010101011111000000000000100";
         f_reg(109) <= "00000000101011100000100000100000";
         f_reg(110) <= "00000010011111000111100000100000";
         f_reg(111) <= "00000001010000100011100000100000";
         f_reg(112) <= "00000011000100001010100000100000";
         f_reg(113) <= "00000000000000000000000000000000";
         f_reg(114) <= "00000000000000000000000000000000";
         f_reg(115) <= "00100000100001011000110010110101";
         f_reg(116) <= "00100010010100111000110010110101";
         f_reg(117) <= "00000000000000000000000000000000";
         f_reg(118) <= "00000000000000000000000000000000";
         f_reg(119) <= "00000000110010110111000000100010";
         f_reg(120) <= "00000010100110011110000000100010";
         f_reg(121) <= "00000001100000000101000000100110";
         f_reg(122) <= "00000011010000001100000000100110";
         f_reg(123) <= "00100100001000100110000001100110";
         f_reg(124) <= "00100101111100000110000001100110";
         f_reg(125) <= "00010101001101110000000011001000";
         f_reg(126) <= "10101100000010010000001100101100";
         f_reg(127) <= "00110000001001001011001011011010";
         f_reg(128) <= "00110001111100101011001011011010";
         f_reg(129) <= "00000000000000000000000000000000";
         f_reg(130) <= "00000000000000000000000000000000";
         f_reg(131) <= "00010101010110000000000011000010";
         f_reg(132) <= "10101100000010100000001100110000";
         f_reg(133) <= "00010101110111000000000011000000";
         f_reg(134) <= "10101100000011100000001100110100";
         f_reg(135) <= "00100100101001101010000010110001";
         f_reg(136) <= "00100110011101001010000010110001";
         f_reg(137) <= "00010100100100100000000010111100";
         f_reg(138) <= "10101100000001000000001100111000";
         f_reg(139) <= "00000000000000000000000000000000";
         f_reg(140) <= "00000000000000000000000000000000";
         f_reg(141) <= "00000000110010000101100000000110";
         f_reg(142) <= "00000010100101101100100000000110";
         f_reg(143) <= "00111100000010011101000111110000";
         f_reg(144) <= "00111100000101111101000111110000";
         f_reg(145) <= "00010101011110010000000010110100";
         f_reg(146) <= "10101100000010110000001100111100";
         f_reg(147) <= "00101000011000011011011110100110";
         f_reg(148) <= "00101010001011111011011110100110";
         f_reg(149) <= "00101000101011101010010111101111";
         f_reg(150) <= "00101010011111001010010111101111";
         f_reg(151) <= "00010101110111000000000010101110";
         f_reg(152) <= "10101100000011100000001101000000";
         f_reg(153) <= "00111100000001000111001101000100";
         f_reg(154) <= "00111100000100100111001101000100";
         f_reg(155) <= "00000001010010010011000000100011";
         f_reg(156) <= "00000011000101111010000000100011";
         f_reg(157) <= "00000000000000000000000000000000";
         f_reg(158) <= "00000000000000000000000000000000";
         f_reg(159) <= "00000000010011000101100000000110";
         f_reg(160) <= "00000010000110101100100000000110";
         f_reg(161) <= "00010101000101100000000010100100";
         f_reg(162) <= "10101100000010000000001101000100";
         f_reg(163) <= "00000001011001110001100000100111";
         f_reg(164) <= "00000011001101011000100000100111";
         f_reg(165) <= "00010100111101010000000010100000";
         f_reg(166) <= "10101100000001110000001101001000";
         f_reg(167) <= "00010100011100010000000010011110";
         f_reg(168) <= "10101100000000110000001101001100";
         f_reg(169) <= "00000000100011010010100000101010";
         f_reg(170) <= "00000010010110111001100000101010";
         f_reg(171) <= "00000000110000010011000000100001";
         f_reg(172) <= "00000010100011111010000000100001";
         f_reg(173) <= "00010101000101100000000010011000";
         f_reg(174) <= "10101100000010000000001101010000";
         f_reg(175) <= "00000000000000000000000000000000";
         f_reg(176) <= "00000000000000000000000000000000";
         f_reg(177) <= "00000000000000000000000000000000";
         f_reg(178) <= "00000000000000000000000000000000";
         f_reg(179) <= "00000000000001010111000011000000";
         f_reg(180) <= "00000000000100111110000011000000";
         f_reg(181) <= "00000000000001010101001001000011";
         f_reg(182) <= "00000000000100111100001001000011";
         f_reg(183) <= "00100000110010011100101101101010";
         f_reg(184) <= "00100010100101111100101101101010";
         f_reg(185) <= "00010101110111000000000010001100";
         f_reg(186) <= "10101100000011100000001101010100";
         f_reg(187) <= "00010101010110000000000010001010";
         f_reg(188) <= "10101100000010100000001101011000";
         f_reg(189) <= "00010101001101110000000010001000";
         f_reg(190) <= "10101100000010010000001101011100";
         f_reg(191) <= "00010100110101000000000010000110";
         f_reg(192) <= "10101100000001100000001101100000";
         f_reg(193) <= "00100011110111011111111100000110";
         f_reg(194) <= "00010011101000000000000000011000";
         f_reg(195) <= "00100011110111011111111000001100";
         f_reg(196) <= "00010011101000000000000000010110";
         f_reg(197) <= "00100011110111011111110100010010";
         f_reg(198) <= "00010011101000000000000000010100";
         f_reg(199) <= "00100011110111101111111111111111";
         f_reg(200) <= "00100011111111111111111111111111";
         f_reg(201) <= "00010111110111110000000001111100";
         f_reg(202) <= "00011111111000001111111101111101";
         f_reg(203) <= "00010000000000000000000100000111";
         f_reg(204) <= "00000000000000000000000000000000";
         f_reg(205) <= "00000000000000000000000000000000";
         f_reg(206) <= "00000000000000000000000000000000";
         f_reg(207) <= "00000000000000000000000000000000";
         f_reg(208) <= "00000000000000000000000000000000";
         f_reg(209) <= "00000000000000000000000000000000";
         f_reg(210) <= "00000000000000000000000000000000";
         f_reg(211) <= "00000000000000000000000000000000";
         f_reg(212) <= "00000000000000000000000000000000";
         f_reg(213) <= "00000000000000000000000000000000";
         f_reg(214) <= "00000000000000000000000000000000";
         f_reg(215) <= "00000000000000000000000000000000";
         f_reg(216) <= "00000000000000000000000000000000";
         f_reg(217) <= "00000000000000000000000000000000";
         f_reg(218) <= "10001100000111010000011010111000";
         f_reg(219) <= "00011111101000000000000000000011";
         f_reg(220) <= "00100000000111010000000000111100";
         f_reg(221) <= "00010000000000000000000000000010";
         f_reg(222) <= "00100000000111010000000000000000";
         f_reg(223) <= "00010100001011110000000001100110";
         f_reg(224) <= "10101111101000010000011001000000";
         f_reg(225) <= "10001100000111010000011010111000";
         f_reg(226) <= "00011111101000000000000000000011";
         f_reg(227) <= "00100000000111010000000000111100";
         f_reg(228) <= "00010000000000000000000000000010";
         f_reg(229) <= "00100000000111010000000000000000";
         f_reg(230) <= "00010100010100000000000001011111";
         f_reg(231) <= "10101111101000100000011001000100";
         f_reg(232) <= "10001100000111010000011010111000";
         f_reg(233) <= "00011111101000000000000000000011";
         f_reg(234) <= "00100000000111010000000000111100";
         f_reg(235) <= "00010000000000000000000000000010";
         f_reg(236) <= "00100000000111010000000000000000";
         f_reg(237) <= "00010100011100010000000001011000";
         f_reg(238) <= "10101111101000110000011001001000";
         f_reg(239) <= "10001100000111010000011010111000";
         f_reg(240) <= "00011111101000000000000000000011";
         f_reg(241) <= "00100000000111010000000000111100";
         f_reg(242) <= "00010000000000000000000000000010";
         f_reg(243) <= "00100000000111010000000000000000";
         f_reg(244) <= "00010100100100100000000001010001";
         f_reg(245) <= "10101111101001000000011001001100";
         f_reg(246) <= "10001100000111010000011010111000";
         f_reg(247) <= "00011111101000000000000000000011";
         f_reg(248) <= "00100000000111010000000000111100";
         f_reg(249) <= "00010000000000000000000000000010";
         f_reg(250) <= "00100000000111010000000000000000";
         f_reg(251) <= "00010100101100110000000001001010";
         f_reg(252) <= "10101111101001010000011001010000";
         f_reg(253) <= "10001100000111010000011010111000";
         f_reg(254) <= "00011111101000000000000000000011";
         f_reg(255) <= "00100000000111010000000000111100";
         f_reg(256) <= "00010000000000000000000000000010";
         f_reg(257) <= "00100000000111010000000000000000";
         f_reg(258) <= "00010100110101000000000001000011";
         f_reg(259) <= "10101111101001100000011001010100";
         f_reg(260) <= "10001100000111010000011010111000";
         f_reg(261) <= "00011111101000000000000000000011";
         f_reg(262) <= "00100000000111010000000000111100";
         f_reg(263) <= "00010000000000000000000000000010";
         f_reg(264) <= "00100000000111010000000000000000";
         f_reg(265) <= "00010100111101010000000000111100";
         f_reg(266) <= "10101111101001110000011001011000";
         f_reg(267) <= "10001100000111010000011010111000";
         f_reg(268) <= "00011111101000000000000000000011";
         f_reg(269) <= "00100000000111010000000000111100";
         f_reg(270) <= "00010000000000000000000000000010";
         f_reg(271) <= "00100000000111010000000000000000";
         f_reg(272) <= "00010101000101100000000000110101";
         f_reg(273) <= "10101111101010000000011001011100";
         f_reg(274) <= "10001100000111010000011010111000";
         f_reg(275) <= "00011111101000000000000000000011";
         f_reg(276) <= "00100000000111010000000000111100";
         f_reg(277) <= "00010000000000000000000000000010";
         f_reg(278) <= "00100000000111010000000000000000";
         f_reg(279) <= "00010101001101110000000000101110";
         f_reg(280) <= "10101111101010010000011001100000";
         f_reg(281) <= "10001100000111010000011010111000";
         f_reg(282) <= "00011111101000000000000000000011";
         f_reg(283) <= "00100000000111010000000000111100";
         f_reg(284) <= "00010000000000000000000000000010";
         f_reg(285) <= "00100000000111010000000000000000";
         f_reg(286) <= "00010101010110000000000000100111";
         f_reg(287) <= "10101111101010100000011001100100";
         f_reg(288) <= "10001100000111010000011010111000";
         f_reg(289) <= "00011111101000000000000000000011";
         f_reg(290) <= "00100000000111010000000000111100";
         f_reg(291) <= "00010000000000000000000000000010";
         f_reg(292) <= "00100000000111010000000000000000";
         f_reg(293) <= "00010101011110010000000000100000";
         f_reg(294) <= "10101111101010110000011001101000";
         f_reg(295) <= "10001100000111010000011010111000";
         f_reg(296) <= "00011111101000000000000000000011";
         f_reg(297) <= "00100000000111010000000000111100";
         f_reg(298) <= "00010000000000000000000000000010";
         f_reg(299) <= "00100000000111010000000000000000";
         f_reg(300) <= "00010101100110100000000000011001";
         f_reg(301) <= "10101111101011000000011001101100";
         f_reg(302) <= "10001100000111010000011010111000";
         f_reg(303) <= "00011111101000000000000000000011";
         f_reg(304) <= "00100000000111010000000000111100";
         f_reg(305) <= "00010000000000000000000000000010";
         f_reg(306) <= "00100000000111010000000000000000";
         f_reg(307) <= "00010101101110110000000000010010";
         f_reg(308) <= "10101111101011010000011001110000";
         f_reg(309) <= "10001100000111010000011010111000";
         f_reg(310) <= "00011111101000000000000000000011";
         f_reg(311) <= "00100000000111010000000000111100";
         f_reg(312) <= "00010000000000000000000000000010";
         f_reg(313) <= "00100000000111010000000000000000";
         f_reg(314) <= "00010101110111000000000000001011";
         f_reg(315) <= "10101111101011100000011001110100";
         f_reg(316) <= "10001100000111010000011010111000";
         f_reg(317) <= "00011111101000000000000000000011";
         f_reg(318) <= "00100000000111010000000000111100";
         f_reg(319) <= "00010000000000000000000000000010";
         f_reg(320) <= "00100000000111010000000000000000";
         f_reg(321) <= "00010111110111110000000000000100";
         f_reg(322) <= "10101111101111100000011001111000";
         f_reg(323) <= "10101100000111010000011010111000";
         f_reg(324) <= "00010000000000001111111110000011";
         f_reg(325) <= "10001100000111010000011010111000";
         f_reg(326) <= "10001111101000010000011001000000";
         f_reg(327) <= "10001100000111010000011010111000";
         f_reg(328) <= "10001111101011110000011001000000";
         f_reg(329) <= "00010100001011111111111111111100";
         f_reg(330) <= "10001100000111010000011010111000";
         f_reg(331) <= "10001111101000100000011001000100";
         f_reg(332) <= "10001100000111010000011010111000";
         f_reg(333) <= "10001111101100000000011001000100";
         f_reg(334) <= "00010100010100001111111111111100";
         f_reg(335) <= "10001100000111010000011010111000";
         f_reg(336) <= "10001111101000110000011001001000";
         f_reg(337) <= "10001100000111010000011010111000";
         f_reg(338) <= "10001111101100010000011001001000";
         f_reg(339) <= "00010100011100011111111111111100";
         f_reg(340) <= "10001100000111010000011010111000";
         f_reg(341) <= "10001111101001000000011001001100";
         f_reg(342) <= "10001100000111010000011010111000";
         f_reg(343) <= "10001111101100100000011001001100";
         f_reg(344) <= "00010100100100101111111111111100";
         f_reg(345) <= "10001100000111010000011010111000";
         f_reg(346) <= "10001111101001010000011001010000";
         f_reg(347) <= "10001100000111010000011010111000";
         f_reg(348) <= "10001111101100110000011001010000";
         f_reg(349) <= "00010100101100111111111111111100";
         f_reg(350) <= "10001100000111010000011010111000";
         f_reg(351) <= "10001111101001100000011001010100";
         f_reg(352) <= "10001100000111010000011010111000";
         f_reg(353) <= "10001111101101000000011001010100";
         f_reg(354) <= "00010100110101001111111111111100";
         f_reg(355) <= "10001100000111010000011010111000";
         f_reg(356) <= "10001111101001110000011001011000";
         f_reg(357) <= "10001100000111010000011010111000";
         f_reg(358) <= "10001111101101010000011001011000";
         f_reg(359) <= "00010100111101011111111111111100";
         f_reg(360) <= "10001100000111010000011010111000";
         f_reg(361) <= "10001111101010000000011001011100";
         f_reg(362) <= "10001100000111010000011010111000";
         f_reg(363) <= "10001111101101100000011001011100";
         f_reg(364) <= "00010101000101101111111111111100";
         f_reg(365) <= "10001100000111010000011010111000";
         f_reg(366) <= "10001111101010010000011001100000";
         f_reg(367) <= "10001100000111010000011010111000";
         f_reg(368) <= "10001111101101110000011001100000";
         f_reg(369) <= "00010101001101111111111111111100";
         f_reg(370) <= "10001100000111010000011010111000";
         f_reg(371) <= "10001111101010100000011001100100";
         f_reg(372) <= "10001100000111010000011010111000";
         f_reg(373) <= "10001111101110000000011001100100";
         f_reg(374) <= "00010101010110001111111111111100";
         f_reg(375) <= "10001100000111010000011010111000";
         f_reg(376) <= "10001111101010110000011001101000";
         f_reg(377) <= "10001100000111010000011010111000";
         f_reg(378) <= "10001111101110010000011001101000";
         f_reg(379) <= "00010101011110011111111111111100";
         f_reg(380) <= "10001100000111010000011010111000";
         f_reg(381) <= "10001111101011000000011001101100";
         f_reg(382) <= "10001100000111010000011010111000";
         f_reg(383) <= "10001111101110100000011001101100";
         f_reg(384) <= "00010101100110101111111111111100";
         f_reg(385) <= "10001100000111010000011010111000";
         f_reg(386) <= "10001111101011010000011001110000";
         f_reg(387) <= "10001100000111010000011010111000";
         f_reg(388) <= "10001111101110110000011001110000";
         f_reg(389) <= "00010101101110111111111111111100";
         f_reg(390) <= "10001100000111010000011010111000";
         f_reg(391) <= "10001111101011100000011001110100";
         f_reg(392) <= "10001100000111010000011010111000";
         f_reg(393) <= "10001111101111000000011001110100";
         f_reg(394) <= "00010101110111001111111111111100";
         f_reg(395) <= "10001100000111010000011010111000";
         f_reg(396) <= "10001111101111100000011001111000";
         f_reg(397) <= "10001100000111010000011010111000";
         f_reg(398) <= "10001111101111110000011001111000";
         f_reg(399) <= "00010111110111111111111111111100";
         f_reg(400) <= "00010000000000001111111100110111";
         f_reg(401) <= "00000000000000000000000000000000";
         f_reg(402) <= "00000000000000000000000000000000";
         f_reg(403) <= "00000000000000000000000000000000";
         f_reg(404) <= "00000000000000000000000000000000";
         f_reg(405) <= "00000000000000000000000000000000";
         f_reg(406) <= "00000000000000000000000000000000";
         f_reg(407) <= "00000000000000000000000000000000";
         f_reg(408) <= "00000000000000000000000000000000";
         f_reg(409) <= "00000000000000000000000000000000";
         f_reg(410) <= "00000000000000000000000000000000";
         f_reg(411) <= "00000000000000000000000000000000";
         f_reg(412) <= "00000000000000000000000000000000";
         f_reg(413) <= "00000000000000000000000000000000";
         f_reg(414) <= "00000000000000000000000000000000";
         f_reg(415) <= "00000000000000000000000000000000";
         f_reg(416) <= "00000000000000000000000000000000";
         f_reg(417) <= "00000000000000000000000000000000";
         f_reg(418) <= "00000000000000000000000000000000";
         f_reg(419) <= "00000000000000000000000000000000";
         f_reg(420) <= "00000000000000000000000000000000";
         f_reg(421) <= "00000000000000000000000000000000";
         f_reg(422) <= "00000000000000000000000000000000";
         f_reg(423) <= "00000000000000000000000000000000";
         f_reg(424) <= "00000000000000000000000000000000";
         f_reg(425) <= "00000000000000000000000000000000";
         f_reg(426) <= "00000000000000000000000000000000";
         f_reg(427) <= "00000000000000000000000000000000";
         f_reg(428) <= "00000000000000000000000000000000";
         f_reg(429) <= "00000000000000000000000000000000";
         f_reg(430) <= "00000000000000000000000000000000";
         f_reg(431) <= "00000000000000000000001111100111";
         f_reg(432) <= "00000000000000000000000000000000";
         f_reg(433) <= "00000000000000000000000000000000";
         f_reg(434) <= "00000000000000000000000000000000";
         f_reg(435) <= "00000000000000000000000000000000";
         f_reg(436) <= "00000000000000000000000000000000";
         f_reg(437) <= "00000000000000000000000000000000";
         f_reg(438) <= "00000000000000000000000000000000";
         f_reg(439) <= "00000000000000000000000000000000";
         f_reg(440) <= "00000000000000000000000000000000";
         f_reg(441) <= "00000000000000000000000000000000";
         f_reg(442) <= "00000000000000000000000000000000";
         f_reg(443) <= "00000000000000000000000000000000";
         f_reg(444) <= "00000000000000000000000000000000";
         f_reg(445) <= "00000000000000000000000000000000";
         f_reg(446) <= "00000000000000000000000000000000";
         f_reg(447) <= "00000000000000000000000000000000";
         f_reg(448) <= "00000000000000000000000000000000";
         f_reg(449) <= "00000000000000000000000000000000";
         f_reg(450) <= "00000000000000000000000000000000";
         f_reg(451) <= "00000000000000000000000000000000";
         f_reg(452) <= "00000000000000000000000000000000";
         f_reg(453) <= "00000000000000000000000000000000";
         f_reg(454) <= "00000000000000000000000000000000";
         f_reg(455) <= "00000000000000000000000000000000";
         f_reg(456) <= "00000000000000000000000000000000";
         f_reg(457) <= "00000000000000000000000000000000";
         f_reg(458) <= "00000000000000000000000000000000";
         f_reg(459) <= "00000000000000000000000000000000";
         f_reg(460) <= "00000000000000000000000000000000";
         f_reg(461) <= "00000000000000000000000000000000";
         f_reg(462) <= "00000000000000000000000000000000";
         f_reg(463) <= "00000000000000000000000000000000";
         f_reg(464) <= "00000000000000000000000000000000";
         f_reg(465) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 -31521
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SLTI R2 R0 5593
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SLTIU R3 R0 2299
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SLLV R4 R0 R2
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SUBU R5 R2 R0
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- ADD R6 R2 R5
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- SLT R7 R4 R4
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- ADDU R8 R7 R4
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- SLTIU R9 R0 -17025
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- NOR R10 R8 R0
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- AND R11 R10 R9
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- ADDIU R12 R7 27880
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- ADDI R13 R5 32229
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- SLTI R14 R6 4484
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- ORI R15 R5 21919
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- OR R16 R8 R8
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SUB R17 R8 R0
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- ADDU R18 R15 R13
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SLLV R19 R1 R7
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- ADD R20 R5 R14
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- ADD R21 R16 R19
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- NOP
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- ADDI R22 R4 -29515
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- NOP
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- SUB R23 R18 R11
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- XOR R24 R12 R0
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- ADDIU R25 R20 24678
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- SW R17 R0 812
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- ANDI R26 R20 -19750
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- NOP
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- SW R24 R0 816
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- SW R23 R0 820
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- ADDIU R27 R22 -24399
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- SW R26 R0 824
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- NOP
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- SRLV R28 R8 R27
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- LUI R29 -11792
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- SW R28 R0 828
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- SLTI R30 R3 -18522
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- SLTI R2 R22 -23057
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SW R2 R0 832
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- LUI R10 29508
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- SUBU R9 R24 R29
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- NOP
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- SRLV R6 R12 R25
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- SW R8 R0 836
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- NOR R15 R6 R21
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- SW R21 R0 840
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SW R15 R0 844
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- SLT R1 R10 R13
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- ADDU R9 R9 R30
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SW R8 R0 848
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- NOP
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- NOP
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SLL R7 R1 3
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- SRA R5 R1 9
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- ADDI R14 R9 -13462
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SW R7 R0 852
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- SW R5 R0 856
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- SW R14 R0 860
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- SW R9 R0 864
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- BGTZ R31 -62
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- BEQ R0 R0 400
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- LUI R30 999
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- LUI R31 999
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- LUI R1 -31521
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- LUI R15 -31521
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SLTI R2 R0 5593
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- SLTI R16 R0 5593
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- SLTIU R3 R0 2299
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- SLTIU R17 R0 2299
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- SLLV R4 R0 R2
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- SLLV R18 R0 R16
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- SUBU R5 R2 R0
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- SUBU R19 R16 R0
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- ADD R6 R2 R5
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- ADD R20 R16 R19
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SLT R7 R4 R4
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- SLT R21 R18 R18
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- ADDU R8 R7 R4
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- ADDU R22 R21 R18
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SLTIU R9 R0 -17025
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- SLTIU R23 R0 -17025
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- NOR R10 R8 R0
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- NOR R24 R22 R0
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- AND R11 R10 R9
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- AND R25 R24 R23
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- ADDIU R12 R7 27880
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- ADDIU R26 R21 27880
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- ADDI R13 R5 32229
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- ADDI R27 R19 32229
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SLTI R14 R6 4484
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SLTI R28 R20 4484
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- ORI R2 R5 21919
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- ORI R16 R19 21919
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- OR R10 R8 R8
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- OR R24 R22 R22
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SUB R9 R8 R0
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- SUB R23 R22 R0
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- ADDU R6 R2 R13
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- ADDU R20 R16 R27
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- SLLV R2 R1 R7
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- SLLV R16 R15 R21
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- ADD R1 R5 R14
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- ADD R15 R19 R28
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- ADD R7 R10 R2
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- ADD R21 R24 R16
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- NOP
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- NOP
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- ADDI R5 R4 -29515
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- ADDI R19 R18 -29515
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- NOP
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- NOP
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- SUB R14 R6 R11
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- SUB R28 R20 R25
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- XOR R10 R12 R0
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- XOR R24 R26 R0
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- ADDIU R2 R1 24678
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- ADDIU R16 R15 24678
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- BNE R9 R23 200
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- SW R9 R0 812
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- ANDI R4 R1 -19750
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- ANDI R18 R15 -19750
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- NOP
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- NOP
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- BNE R10 R24 194
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- SW R10 R0 816
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- BNE R14 R28 192
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- SW R14 R0 820
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- ADDIU R6 R5 -24399
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- ADDIU R20 R19 -24399
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- BNE R4 R18 188
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SW R4 R0 824
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- NOP
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- NOP
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- SRLV R11 R8 R6
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- SRLV R25 R22 R20
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- LUI R9 -11792
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- LUI R23 -11792
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- BNE R11 R25 180
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- SW R11 R0 828
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- SLTI R1 R3 -18522
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- SLTI R15 R17 -18522
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- SLTI R14 R5 -23057
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- SLTI R28 R19 -23057
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- BNE R14 R28 174
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- SW R14 R0 832
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- LUI R4 29508
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- LUI R18 29508
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- SUBU R6 R10 R9
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- SUBU R20 R24 R23
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- NOP
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- NOP
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- SRLV R11 R12 R2
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- SRLV R25 R26 R16
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- BNE R8 R22 164
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- SW R8 R0 836
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- NOR R3 R11 R7
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- NOR R17 R25 R21
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- BNE R7 R21 160
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- SW R7 R0 840
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- BNE R3 R17 158
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- SW R3 R0 844
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- SLT R5 R4 R13
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- SLT R19 R18 R27
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- ADDU R6 R6 R1
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- ADDU R20 R20 R15
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- BNE R8 R22 152
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- SW R8 R0 848
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- NOP
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- NOP
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- NOP
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- NOP
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- SLL R14 R5 3
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- SLL R28 R19 3
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- SRA R10 R5 9
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SRA R24 R19 9
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- ADDI R9 R6 -13462
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- ADDI R23 R20 -13462
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- BNE R14 R28 140
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- SW R14 R0 852
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- BNE R10 R24 138
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- SW R10 R0 856
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- BNE R9 R23 136
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- SW R9 R0 860
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- BNE R6 R20 134
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- SW R6 R0 864
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- BEQ R29 R0 24
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- BEQ R29 R0 22
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- BEQ R29 R0 20
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- BNE R30 R31 124
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- BGTZ R31 -131
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- BEQ R0 R0 263
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- NOP
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- NOP
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- NOP
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- NOP
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- NOP
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- NOP
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- NOP
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- NOP
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- NOP
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- NOP
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- NOP
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- NOP
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- NOP
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- NOP
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- SW R1 R29 1600
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- SW R2 R29 1604
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- SW R3 R29 1608
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- SW R4 R29 1612
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- SW R5 R29 1616
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- SW R6 R29 1620
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- SW R7 R29 1624
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- SW R8 R29 1628
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- SW R9 R29 1632
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- SW R10 R29 1636
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- SW R11 R29 1640
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- SW R12 R29 1644
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- SW R13 R29 1648
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- SW R14 R29 1652
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- SW R30 R29 1656
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- SW R29 R0 1720
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- BEQ R0 R0 -125
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- LW R1 R29 1600
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- LW R15 R29 1600
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- LW R2 R29 1604
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- LW R16 R29 1604
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- LW R3 R29 1608
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- LW R17 R29 1608
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- LW R4 R29 1612
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- LW R18 R29 1612
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- LW R5 R29 1616
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- LW R19 R29 1616
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- LW R6 R29 1620
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- LW R20 R29 1620
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- LW R7 R29 1624
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- LW R21 R29 1624
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- LW R8 R29 1628
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- LW R22 R29 1628
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- LW R9 R29 1632
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- LW R23 R29 1632
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- LW R10 R29 1636
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- LW R24 R29 1636
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- LW R11 R29 1640
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- LW R25 R29 1640
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- LW R12 R29 1644
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- LW R26 R29 1644
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- LW R13 R29 1648
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- LW R27 R29 1648
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- LW R14 R29 1652
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- LW R28 R29 1652
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- LW R30 R29 1656
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- LW R29 R0 1720
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- LW R31 R29 1656
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- BEQ R0 R0 -201
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- NOP
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- NOP
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- NOP
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- NOP
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- NOP
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- NOP
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- NOP
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- NOP
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- NOP
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- NOP
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- NOP
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- NOP
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- NOP
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- NOP
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- NOP
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- NOP
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- NOP
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- NOP
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- NOP
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- NOP
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- NOP
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- NOP
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- NOP
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- NOP
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- NOP
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- NOP
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- NOP
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- NOP
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- NOP
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- NOP
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- NOP
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- NOP
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- NOP
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- NOP
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- NOP
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- NOP
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- NOP
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- NOP
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- NOP
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- NOP
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- NOP
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- NOP
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- NOP
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- NOP
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- NOP
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- NOP
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- NOP
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- NOP
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- NOP
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- NOP
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- NOP
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- NOP
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- NOP
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- NOP
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- NOP
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- NOP
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- NOP
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- NOP
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- NOP
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- NOP
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- NOP
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- NOP
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- NOP
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- NOP
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- NOP
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011000010011011111";
                        f_reg(4) <= "00101000000000100001010111011001";
                        f_reg(5) <= "00101100000000110000100011111011";
                        f_reg(6) <= "00000000010000000010000000000100";
                        f_reg(7) <= "00000000010000000010100000100011";
                        f_reg(8) <= "00000000010001010011000000100000";
                        f_reg(9) <= "00000000100001000011100000101010";
                        f_reg(10) <= "00000000111001000100000000100001";
                        f_reg(11) <= "00101100000010011011110101111111";
                        f_reg(12) <= "00000001000000000101000000100111";
                        f_reg(13) <= "00000001010010010101100000100100";
                        f_reg(14) <= "00100100111011000110110011101000";
                        f_reg(15) <= "00100000101011010111110111100101";
                        f_reg(16) <= "00101000110011100001000110000100";
                        f_reg(17) <= "00110100101011110101010110011111";
                        f_reg(18) <= "00000001000010001000000000100101";
                        f_reg(19) <= "00000001000000001000100000100010";
                        f_reg(20) <= "00000001111011011001000000100001";
                        f_reg(21) <= "00000000111000011001100000000100";
                        f_reg(22) <= "00000000101011101010000000100000";
                        f_reg(23) <= "00000010000100111010100000100000";
                        f_reg(24) <= "00000000000000000000000000000000";
                        f_reg(25) <= "00100000100101101000110010110101";
                        f_reg(26) <= "00000000000000000000000000000000";
                        f_reg(27) <= "00000010010010111011100000100010";
                        f_reg(28) <= "00000001100000001100000000100110";
                        f_reg(29) <= "00100110100110010110000001100110";
                        f_reg(30) <= "10101100000100010000001100101100";
                        f_reg(31) <= "00110010100110101011001011011010";
                        f_reg(32) <= "00000000000000000000000000000000";
                        f_reg(33) <= "10101100000110000000001100110000";
                        f_reg(34) <= "10101100000101110000001100110100";
                        f_reg(35) <= "00100110110110111010000010110001";
                        f_reg(36) <= "10101100000110100000001100111000";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00000011011010001110000000000110";
                        f_reg(39) <= "00111100000111011101000111110000";
                        f_reg(40) <= "10101100000111000000001100111100";
                        f_reg(41) <= "00101000011111101011011110100110";
                        f_reg(42) <= "00101010110000101010010111101111";
                        f_reg(43) <= "10101100000000100000001101000000";
                        f_reg(44) <= "00111100000010100111001101000100";
                        f_reg(45) <= "00000011000111010100100000100011";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00000011001011000011000000000110";
                        f_reg(48) <= "10101100000010000000001101000100";
                        f_reg(49) <= "00000000110101010111100000100111";
                        f_reg(50) <= "10101100000101010000001101001000";
                        f_reg(51) <= "10101100000011110000001101001100";
                        f_reg(52) <= "00000001010011010000100000101010";
                        f_reg(53) <= "00000001001111100100100000100001";
                        f_reg(54) <= "10101100000010000000001101010000";
                        f_reg(55) <= "00000000000000000000000000000000";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000010011100011000000";
                        f_reg(58) <= "00000000000000010010101001000011";
                        f_reg(59) <= "00100001001011101100101101101010";
                        f_reg(60) <= "10101100000001110000001101010100";
                        f_reg(61) <= "10101100000001010000001101011000";
                        f_reg(62) <= "10101100000011100000001101011100";
                        f_reg(63) <= "10101100000010010000001101100000";
                        f_reg(64) <= "00100011111111111111111111111111";
                        f_reg(65) <= "00011111111000001111111111000010";
                        f_reg(66) <= "00010000000000000000000110010000";
                        f_reg(67) <= "00111100000111100000001111100111";
                        f_reg(68) <= "00111100000111110000001111100111";
                        f_reg(69) <= "00000000000111101111010000000010";
                        f_reg(70) <= "00000000000111111111110000000010";
                        f_reg(71) <= "00111100000000011000010011011111";
                        f_reg(72) <= "00111100000011111000010011011111";
                        f_reg(73) <= "00101000000000100001010111011001";
                        f_reg(74) <= "00101000000100000001010111011001";
                        f_reg(75) <= "00101100000000110000100011111011";
                        f_reg(76) <= "00101100000100010000100011111011";
                        f_reg(77) <= "00000000010000000010000000000100";
                        f_reg(78) <= "00000010000000001001000000000100";
                        f_reg(79) <= "00000000010000000010100000100011";
                        f_reg(80) <= "00000010000000001001100000100011";
                        f_reg(81) <= "00000000010001010011000000100000";
                        f_reg(82) <= "00000010000100111010000000100000";
                        f_reg(83) <= "00000000100001000011100000101010";
                        f_reg(84) <= "00000010010100101010100000101010";
                        f_reg(85) <= "00000000111001000100000000100001";
                        f_reg(86) <= "00000010101100101011000000100001";
                        f_reg(87) <= "00101100000010011011110101111111";
                        f_reg(88) <= "00101100000101111011110101111111";
                        f_reg(89) <= "00000001000000000101000000100111";
                        f_reg(90) <= "00000010110000001100000000100111";
                        f_reg(91) <= "00000001010010010101100000100100";
                        f_reg(92) <= "00000011000101111100100000100100";
                        f_reg(93) <= "00100100111011000110110011101000";
                        f_reg(94) <= "00100110101110100110110011101000";
                        f_reg(95) <= "00100000101011010111110111100101";
                        f_reg(96) <= "00100010011110110111110111100101";
                        f_reg(97) <= "00101000110011100001000110000100";
                        f_reg(98) <= "00101010100111000001000110000100";
                        f_reg(99) <= "00110100101000100101010110011111";
                        f_reg(100) <= "00110110011100000101010110011111";
                        f_reg(101) <= "00000001000010000101000000100101";
                        f_reg(102) <= "00000010110101101100000000100101";
                        f_reg(103) <= "00000001000000000100100000100010";
                        f_reg(104) <= "00000010110000001011100000100010";
                        f_reg(105) <= "00000000010011010011000000100001";
                        f_reg(106) <= "00000010000110111010000000100001";
                        f_reg(107) <= "00000000111000010001000000000100";
                        f_reg(108) <= "00000010101011111000000000000100";
                        f_reg(109) <= "00000000101011100000100000100000";
                        f_reg(110) <= "00000010011111000111100000100000";
                        f_reg(111) <= "00000001010000100011100000100000";
                        f_reg(112) <= "00000011000100001010100000100000";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00100000100001011000110010110101";
                        f_reg(116) <= "00100010010100111000110010110101";
                        f_reg(117) <= "00000000000000000000000000000000";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000110010110111000000100010";
                        f_reg(120) <= "00000010100110011110000000100010";
                        f_reg(121) <= "00000001100000000101000000100110";
                        f_reg(122) <= "00000011010000001100000000100110";
                        f_reg(123) <= "00100100001000100110000001100110";
                        f_reg(124) <= "00100101111100000110000001100110";
                        f_reg(125) <= "00010101001101110000000011001000";
                        f_reg(126) <= "10101100000010010000001100101100";
                        f_reg(127) <= "00110000001001001011001011011010";
                        f_reg(128) <= "00110001111100101011001011011010";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010101010110000000000011000010";
                        f_reg(132) <= "10101100000010100000001100110000";
                        f_reg(133) <= "00010101110111000000000011000000";
                        f_reg(134) <= "10101100000011100000001100110100";
                        f_reg(135) <= "00100100101001101010000010110001";
                        f_reg(136) <= "00100110011101001010000010110001";
                        f_reg(137) <= "00010100100100100000000010111100";
                        f_reg(138) <= "10101100000001000000001100111000";
                        f_reg(139) <= "00000000000000000000000000000000";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000110010000101100000000110";
                        f_reg(142) <= "00000010100101101100100000000110";
                        f_reg(143) <= "00111100000010011101000111110000";
                        f_reg(144) <= "00111100000101111101000111110000";
                        f_reg(145) <= "00010101011110010000000010110100";
                        f_reg(146) <= "10101100000010110000001100111100";
                        f_reg(147) <= "00101000011000011011011110100110";
                        f_reg(148) <= "00101010001011111011011110100110";
                        f_reg(149) <= "00101000101011101010010111101111";
                        f_reg(150) <= "00101010011111001010010111101111";
                        f_reg(151) <= "00010101110111000000000010101110";
                        f_reg(152) <= "10101100000011100000001101000000";
                        f_reg(153) <= "00111100000001000111001101000100";
                        f_reg(154) <= "00111100000100100111001101000100";
                        f_reg(155) <= "00000001010010010011000000100011";
                        f_reg(156) <= "00000011000101111010000000100011";
                        f_reg(157) <= "00000000000000000000000000000000";
                        f_reg(158) <= "00000000000000000000000000000000";
                        f_reg(159) <= "00000000010011000101100000000110";
                        f_reg(160) <= "00000010000110101100100000000110";
                        f_reg(161) <= "00010101000101100000000010100100";
                        f_reg(162) <= "10101100000010000000001101000100";
                        f_reg(163) <= "00000001011001110001100000100111";
                        f_reg(164) <= "00000011001101011000100000100111";
                        f_reg(165) <= "00010100111101010000000010100000";
                        f_reg(166) <= "10101100000001110000001101001000";
                        f_reg(167) <= "00010100011100010000000010011110";
                        f_reg(168) <= "10101100000000110000001101001100";
                        f_reg(169) <= "00000000100011010010100000101010";
                        f_reg(170) <= "00000010010110111001100000101010";
                        f_reg(171) <= "00000000110000010011000000100001";
                        f_reg(172) <= "00000010100011111010000000100001";
                        f_reg(173) <= "00010101000101100000000010011000";
                        f_reg(174) <= "10101100000010000000001101010000";
                        f_reg(175) <= "00000000000000000000000000000000";
                        f_reg(176) <= "00000000000000000000000000000000";
                        f_reg(177) <= "00000000000000000000000000000000";
                        f_reg(178) <= "00000000000000000000000000000000";
                        f_reg(179) <= "00000000000001010111000011000000";
                        f_reg(180) <= "00000000000100111110000011000000";
                        f_reg(181) <= "00000000000001010101001001000011";
                        f_reg(182) <= "00000000000100111100001001000011";
                        f_reg(183) <= "00100000110010011100101101101010";
                        f_reg(184) <= "00100010100101111100101101101010";
                        f_reg(185) <= "00010101110111000000000010001100";
                        f_reg(186) <= "10101100000011100000001101010100";
                        f_reg(187) <= "00010101010110000000000010001010";
                        f_reg(188) <= "10101100000010100000001101011000";
                        f_reg(189) <= "00010101001101110000000010001000";
                        f_reg(190) <= "10101100000010010000001101011100";
                        f_reg(191) <= "00010100110101000000000010000110";
                        f_reg(192) <= "10101100000001100000001101100000";
                        f_reg(193) <= "00100011110111011111111100000110";
                        f_reg(194) <= "00010011101000000000000000011000";
                        f_reg(195) <= "00100011110111011111111000001100";
                        f_reg(196) <= "00010011101000000000000000010110";
                        f_reg(197) <= "00100011110111011111110100010010";
                        f_reg(198) <= "00010011101000000000000000010100";
                        f_reg(199) <= "00100011110111101111111111111111";
                        f_reg(200) <= "00100011111111111111111111111111";
                        f_reg(201) <= "00010111110111110000000001111100";
                        f_reg(202) <= "00011111111000001111111101111101";
                        f_reg(203) <= "00010000000000000000000100000111";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000000000000000000000000000000";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00000000000000000000000000000000";
                        f_reg(215) <= "00000000000000000000000000000000";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "10001100000111010000011010111000";
                        f_reg(219) <= "00011111101000000000000000000011";
                        f_reg(220) <= "00100000000111010000000000111100";
                        f_reg(221) <= "00010000000000000000000000000010";
                        f_reg(222) <= "00100000000111010000000000000000";
                        f_reg(223) <= "00010100001011110000000001100110";
                        f_reg(224) <= "10101111101000010000011001000000";
                        f_reg(225) <= "10001100000111010000011010111000";
                        f_reg(226) <= "00011111101000000000000000000011";
                        f_reg(227) <= "00100000000111010000000000111100";
                        f_reg(228) <= "00010000000000000000000000000010";
                        f_reg(229) <= "00100000000111010000000000000000";
                        f_reg(230) <= "00010100010100000000000001011111";
                        f_reg(231) <= "10101111101000100000011001000100";
                        f_reg(232) <= "10001100000111010000011010111000";
                        f_reg(233) <= "00011111101000000000000000000011";
                        f_reg(234) <= "00100000000111010000000000111100";
                        f_reg(235) <= "00010000000000000000000000000010";
                        f_reg(236) <= "00100000000111010000000000000000";
                        f_reg(237) <= "00010100011100010000000001011000";
                        f_reg(238) <= "10101111101000110000011001001000";
                        f_reg(239) <= "10001100000111010000011010111000";
                        f_reg(240) <= "00011111101000000000000000000011";
                        f_reg(241) <= "00100000000111010000000000111100";
                        f_reg(242) <= "00010000000000000000000000000010";
                        f_reg(243) <= "00100000000111010000000000000000";
                        f_reg(244) <= "00010100100100100000000001010001";
                        f_reg(245) <= "10101111101001000000011001001100";
                        f_reg(246) <= "10001100000111010000011010111000";
                        f_reg(247) <= "00011111101000000000000000000011";
                        f_reg(248) <= "00100000000111010000000000111100";
                        f_reg(249) <= "00010000000000000000000000000010";
                        f_reg(250) <= "00100000000111010000000000000000";
                        f_reg(251) <= "00010100101100110000000001001010";
                        f_reg(252) <= "10101111101001010000011001010000";
                        f_reg(253) <= "10001100000111010000011010111000";
                        f_reg(254) <= "00011111101000000000000000000011";
                        f_reg(255) <= "00100000000111010000000000111100";
                        f_reg(256) <= "00010000000000000000000000000010";
                        f_reg(257) <= "00100000000111010000000000000000";
                        f_reg(258) <= "00010100110101000000000001000011";
                        f_reg(259) <= "10101111101001100000011001010100";
                        f_reg(260) <= "10001100000111010000011010111000";
                        f_reg(261) <= "00011111101000000000000000000011";
                        f_reg(262) <= "00100000000111010000000000111100";
                        f_reg(263) <= "00010000000000000000000000000010";
                        f_reg(264) <= "00100000000111010000000000000000";
                        f_reg(265) <= "00010100111101010000000000111100";
                        f_reg(266) <= "10101111101001110000011001011000";
                        f_reg(267) <= "10001100000111010000011010111000";
                        f_reg(268) <= "00011111101000000000000000000011";
                        f_reg(269) <= "00100000000111010000000000111100";
                        f_reg(270) <= "00010000000000000000000000000010";
                        f_reg(271) <= "00100000000111010000000000000000";
                        f_reg(272) <= "00010101000101100000000000110101";
                        f_reg(273) <= "10101111101010000000011001011100";
                        f_reg(274) <= "10001100000111010000011010111000";
                        f_reg(275) <= "00011111101000000000000000000011";
                        f_reg(276) <= "00100000000111010000000000111100";
                        f_reg(277) <= "00010000000000000000000000000010";
                        f_reg(278) <= "00100000000111010000000000000000";
                        f_reg(279) <= "00010101001101110000000000101110";
                        f_reg(280) <= "10101111101010010000011001100000";
                        f_reg(281) <= "10001100000111010000011010111000";
                        f_reg(282) <= "00011111101000000000000000000011";
                        f_reg(283) <= "00100000000111010000000000111100";
                        f_reg(284) <= "00010000000000000000000000000010";
                        f_reg(285) <= "00100000000111010000000000000000";
                        f_reg(286) <= "00010101010110000000000000100111";
                        f_reg(287) <= "10101111101010100000011001100100";
                        f_reg(288) <= "10001100000111010000011010111000";
                        f_reg(289) <= "00011111101000000000000000000011";
                        f_reg(290) <= "00100000000111010000000000111100";
                        f_reg(291) <= "00010000000000000000000000000010";
                        f_reg(292) <= "00100000000111010000000000000000";
                        f_reg(293) <= "00010101011110010000000000100000";
                        f_reg(294) <= "10101111101010110000011001101000";
                        f_reg(295) <= "10001100000111010000011010111000";
                        f_reg(296) <= "00011111101000000000000000000011";
                        f_reg(297) <= "00100000000111010000000000111100";
                        f_reg(298) <= "00010000000000000000000000000010";
                        f_reg(299) <= "00100000000111010000000000000000";
                        f_reg(300) <= "00010101100110100000000000011001";
                        f_reg(301) <= "10101111101011000000011001101100";
                        f_reg(302) <= "10001100000111010000011010111000";
                        f_reg(303) <= "00011111101000000000000000000011";
                        f_reg(304) <= "00100000000111010000000000111100";
                        f_reg(305) <= "00010000000000000000000000000010";
                        f_reg(306) <= "00100000000111010000000000000000";
                        f_reg(307) <= "00010101101110110000000000010010";
                        f_reg(308) <= "10101111101011010000011001110000";
                        f_reg(309) <= "10001100000111010000011010111000";
                        f_reg(310) <= "00011111101000000000000000000011";
                        f_reg(311) <= "00100000000111010000000000111100";
                        f_reg(312) <= "00010000000000000000000000000010";
                        f_reg(313) <= "00100000000111010000000000000000";
                        f_reg(314) <= "00010101110111000000000000001011";
                        f_reg(315) <= "10101111101011100000011001110100";
                        f_reg(316) <= "10001100000111010000011010111000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010111110111110000000000000100";
                        f_reg(322) <= "10101111101111100000011001111000";
                        f_reg(323) <= "10101100000111010000011010111000";
                        f_reg(324) <= "00010000000000001111111110000011";
                        f_reg(325) <= "10001100000111010000011010111000";
                        f_reg(326) <= "10001111101000010000011001000000";
                        f_reg(327) <= "10001100000111010000011010111000";
                        f_reg(328) <= "10001111101011110000011001000000";
                        f_reg(329) <= "00010100001011111111111111111100";
                        f_reg(330) <= "10001100000111010000011010111000";
                        f_reg(331) <= "10001111101000100000011001000100";
                        f_reg(332) <= "10001100000111010000011010111000";
                        f_reg(333) <= "10001111101100000000011001000100";
                        f_reg(334) <= "00010100010100001111111111111100";
                        f_reg(335) <= "10001100000111010000011010111000";
                        f_reg(336) <= "10001111101000110000011001001000";
                        f_reg(337) <= "10001100000111010000011010111000";
                        f_reg(338) <= "10001111101100010000011001001000";
                        f_reg(339) <= "00010100011100011111111111111100";
                        f_reg(340) <= "10001100000111010000011010111000";
                        f_reg(341) <= "10001111101001000000011001001100";
                        f_reg(342) <= "10001100000111010000011010111000";
                        f_reg(343) <= "10001111101100100000011001001100";
                        f_reg(344) <= "00010100100100101111111111111100";
                        f_reg(345) <= "10001100000111010000011010111000";
                        f_reg(346) <= "10001111101001010000011001010000";
                        f_reg(347) <= "10001100000111010000011010111000";
                        f_reg(348) <= "10001111101100110000011001010000";
                        f_reg(349) <= "00010100101100111111111111111100";
                        f_reg(350) <= "10001100000111010000011010111000";
                        f_reg(351) <= "10001111101001100000011001010100";
                        f_reg(352) <= "10001100000111010000011010111000";
                        f_reg(353) <= "10001111101101000000011001010100";
                        f_reg(354) <= "00010100110101001111111111111100";
                        f_reg(355) <= "10001100000111010000011010111000";
                        f_reg(356) <= "10001111101001110000011001011000";
                        f_reg(357) <= "10001100000111010000011010111000";
                        f_reg(358) <= "10001111101101010000011001011000";
                        f_reg(359) <= "00010100111101011111111111111100";
                        f_reg(360) <= "10001100000111010000011010111000";
                        f_reg(361) <= "10001111101010000000011001011100";
                        f_reg(362) <= "10001100000111010000011010111000";
                        f_reg(363) <= "10001111101101100000011001011100";
                        f_reg(364) <= "00010101000101101111111111111100";
                        f_reg(365) <= "10001100000111010000011010111000";
                        f_reg(366) <= "10001111101010010000011001100000";
                        f_reg(367) <= "10001100000111010000011010111000";
                        f_reg(368) <= "10001111101101110000011001100000";
                        f_reg(369) <= "00010101001101111111111111111100";
                        f_reg(370) <= "10001100000111010000011010111000";
                        f_reg(371) <= "10001111101010100000011001100100";
                        f_reg(372) <= "10001100000111010000011010111000";
                        f_reg(373) <= "10001111101110000000011001100100";
                        f_reg(374) <= "00010101010110001111111111111100";
                        f_reg(375) <= "10001100000111010000011010111000";
                        f_reg(376) <= "10001111101010110000011001101000";
                        f_reg(377) <= "10001100000111010000011010111000";
                        f_reg(378) <= "10001111101110010000011001101000";
                        f_reg(379) <= "00010101011110011111111111111100";
                        f_reg(380) <= "10001100000111010000011010111000";
                        f_reg(381) <= "10001111101011000000011001101100";
                        f_reg(382) <= "10001100000111010000011010111000";
                        f_reg(383) <= "10001111101110100000011001101100";
                        f_reg(384) <= "00010101100110101111111111111100";
                        f_reg(385) <= "10001100000111010000011010111000";
                        f_reg(386) <= "10001111101011010000011001110000";
                        f_reg(387) <= "10001100000111010000011010111000";
                        f_reg(388) <= "10001111101110110000011001110000";
                        f_reg(389) <= "00010101101110111111111111111100";
                        f_reg(390) <= "10001100000111010000011010111000";
                        f_reg(391) <= "10001111101011100000011001110100";
                        f_reg(392) <= "10001100000111010000011010111000";
                        f_reg(393) <= "10001111101111000000011001110100";
                        f_reg(394) <= "00010101110111001111111111111100";
                        f_reg(395) <= "10001100000111010000011010111000";
                        f_reg(396) <= "10001111101111100000011001111000";
                        f_reg(397) <= "10001100000111010000011010111000";
                        f_reg(398) <= "10001111101111110000011001111000";
                        f_reg(399) <= "00010111110111111111111111111100";
                        f_reg(400) <= "00010000000000001111111100110111";
                        f_reg(401) <= "00000000000000000000000000000000";
                        f_reg(402) <= "00000000000000000000000000000000";
                        f_reg(403) <= "00000000000000000000000000000000";
                        f_reg(404) <= "00000000000000000000000000000000";
                        f_reg(405) <= "00000000000000000000000000000000";
                        f_reg(406) <= "00000000000000000000000000000000";
                        f_reg(407) <= "00000000000000000000000000000000";
                        f_reg(408) <= "00000000000000000000000000000000";
                        f_reg(409) <= "00000000000000000000000000000000";
                        f_reg(410) <= "00000000000000000000000000000000";
                        f_reg(411) <= "00000000000000000000000000000000";
                        f_reg(412) <= "00000000000000000000000000000000";
                        f_reg(413) <= "00000000000000000000000000000000";
                        f_reg(414) <= "00000000000000000000000000000000";
                        f_reg(415) <= "00000000000000000000000000000000";
                        f_reg(416) <= "00000000000000000000000000000000";
                        f_reg(417) <= "00000000000000000000000000000000";
                        f_reg(418) <= "00000000000000000000000000000000";
                        f_reg(419) <= "00000000000000000000000000000000";
                        f_reg(420) <= "00000000000000000000000000000000";
                        f_reg(421) <= "00000000000000000000000000000000";
                        f_reg(422) <= "00000000000000000000000000000000";
                        f_reg(423) <= "00000000000000000000000000000000";
                        f_reg(424) <= "00000000000000000000000000000000";
                        f_reg(425) <= "00000000000000000000000000000000";
                        f_reg(426) <= "00000000000000000000000000000000";
                        f_reg(427) <= "00000000000000000000000000000000";
                        f_reg(428) <= "00000000000000000000000000000000";
                        f_reg(429) <= "00000000000000000000000000000000";
                        f_reg(430) <= "00000000000000000000000000000000";
                        f_reg(431) <= "00000000000000000000001111100111";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011000010011011111";
                        f_reg(4) <= "00101000000000100001010111011001";
                        f_reg(5) <= "00101100000000110000100011111011";
                        f_reg(6) <= "00000000010000000010000000000100";
                        f_reg(7) <= "00000000010000000010100000100011";
                        f_reg(8) <= "00000000010001010011000000100000";
                        f_reg(9) <= "00000000100001000011100000101010";
                        f_reg(10) <= "00000000111001000100000000100001";
                        f_reg(11) <= "00101100000010011011110101111111";
                        f_reg(12) <= "00000001000000000101000000100111";
                        f_reg(13) <= "00000001010010010101100000100100";
                        f_reg(14) <= "00100100111011000110110011101000";
                        f_reg(15) <= "00100000101011010111110111100101";
                        f_reg(16) <= "00101000110011100001000110000100";
                        f_reg(17) <= "00110100101011110101010110011111";
                        f_reg(18) <= "00000001000010001000000000100101";
                        f_reg(19) <= "00000001000000001000100000100010";
                        f_reg(20) <= "00000001111011011001000000100001";
                        f_reg(21) <= "00000000111000011001100000000100";
                        f_reg(22) <= "00000000101011101010000000100000";
                        f_reg(23) <= "00000010000100111010100000100000";
                        f_reg(24) <= "00000000000000000000000000000000";
                        f_reg(25) <= "00100000100101101000110010110101";
                        f_reg(26) <= "00000000000000000000000000000000";
                        f_reg(27) <= "00000010010010111011100000100010";
                        f_reg(28) <= "00000001100000001100000000100110";
                        f_reg(29) <= "00100110100110010110000001100110";
                        f_reg(30) <= "10101100000100010000001100101100";
                        f_reg(31) <= "00110010100110101011001011011010";
                        f_reg(32) <= "00000000000000000000000000000000";
                        f_reg(33) <= "10101100000110000000001100110000";
                        f_reg(34) <= "10101100000101110000001100110100";
                        f_reg(35) <= "00100110110110111010000010110001";
                        f_reg(36) <= "10101100000110100000001100111000";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00000011011010001110000000000110";
                        f_reg(39) <= "00111100000111011101000111110000";
                        f_reg(40) <= "10101100000111000000001100111100";
                        f_reg(41) <= "00101000011111101011011110100110";
                        f_reg(42) <= "00101010110000101010010111101111";
                        f_reg(43) <= "10101100000000100000001101000000";
                        f_reg(44) <= "00111100000010100111001101000100";
                        f_reg(45) <= "00000011000111010100100000100011";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00000011001011000011000000000110";
                        f_reg(48) <= "10101100000010000000001101000100";
                        f_reg(49) <= "00000000110101010111100000100111";
                        f_reg(50) <= "10101100000101010000001101001000";
                        f_reg(51) <= "10101100000011110000001101001100";
                        f_reg(52) <= "00000001010011010000100000101010";
                        f_reg(53) <= "00000001001111100100100000100001";
                        f_reg(54) <= "10101100000010000000001101010000";
                        f_reg(55) <= "00000000000000000000000000000000";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000010011100011000000";
                        f_reg(58) <= "00000000000000010010101001000011";
                        f_reg(59) <= "00100001001011101100101101101010";
                        f_reg(60) <= "10101100000001110000001101010100";
                        f_reg(61) <= "10101100000001010000001101011000";
                        f_reg(62) <= "10101100000011100000001101011100";
                        f_reg(63) <= "10101100000010010000001101100000";
                        f_reg(64) <= "00100011111111111111111111111111";
                        f_reg(65) <= "00011111111000001111111111000010";
                        f_reg(66) <= "00010000000000000000000110010000";
                        f_reg(67) <= "00111100000111100000001111100111";
                        f_reg(68) <= "00111100000111110000001111100111";
                        f_reg(69) <= "00000000000111101111010000000010";
                        f_reg(70) <= "00000000000111111111110000000010";
                        f_reg(71) <= "00111100000000011000010011011111";
                        f_reg(72) <= "00111100000011111000010011011111";
                        f_reg(73) <= "00101000000000100001010111011001";
                        f_reg(74) <= "00101000000100000001010111011001";
                        f_reg(75) <= "00101100000000110000100011111011";
                        f_reg(76) <= "00101100000100010000100011111011";
                        f_reg(77) <= "00000000010000000010000000000100";
                        f_reg(78) <= "00000010000000001001000000000100";
                        f_reg(79) <= "00000000010000000010100000100011";
                        f_reg(80) <= "00000010000000001001100000100011";
                        f_reg(81) <= "00000000010001010011000000100000";
                        f_reg(82) <= "00000010000100111010000000100000";
                        f_reg(83) <= "00000000100001000011100000101010";
                        f_reg(84) <= "00000010010100101010100000101010";
                        f_reg(85) <= "00000000111001000100000000100001";
                        f_reg(86) <= "00000010101100101011000000100001";
                        f_reg(87) <= "00101100000010011011110101111111";
                        f_reg(88) <= "00101100000101111011110101111111";
                        f_reg(89) <= "00000001000000000101000000100111";
                        f_reg(90) <= "00000010110000001100000000100111";
                        f_reg(91) <= "00000001010010010101100000100100";
                        f_reg(92) <= "00000011000101111100100000100100";
                        f_reg(93) <= "00100100111011000110110011101000";
                        f_reg(94) <= "00100110101110100110110011101000";
                        f_reg(95) <= "00100000101011010111110111100101";
                        f_reg(96) <= "00100010011110110111110111100101";
                        f_reg(97) <= "00101000110011100001000110000100";
                        f_reg(98) <= "00101010100111000001000110000100";
                        f_reg(99) <= "00110100101000100101010110011111";
                        f_reg(100) <= "00110110011100000101010110011111";
                        f_reg(101) <= "00000001000010000101000000100101";
                        f_reg(102) <= "00000010110101101100000000100101";
                        f_reg(103) <= "00000001000000000100100000100010";
                        f_reg(104) <= "00000010110000001011100000100010";
                        f_reg(105) <= "00000000010011010011000000100001";
                        f_reg(106) <= "00000010000110111010000000100001";
                        f_reg(107) <= "00000000111000010001000000000100";
                        f_reg(108) <= "00000010101011111000000000000100";
                        f_reg(109) <= "00000000101011100000100000100000";
                        f_reg(110) <= "00000010011111000111100000100000";
                        f_reg(111) <= "00000001010000100011100000100000";
                        f_reg(112) <= "00000011000100001010100000100000";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00100000100001011000110010110101";
                        f_reg(116) <= "00100010010100111000110010110101";
                        f_reg(117) <= "00000000000000000000000000000000";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000110010110111000000100010";
                        f_reg(120) <= "00000010100110011110000000100010";
                        f_reg(121) <= "00000001100000000101000000100110";
                        f_reg(122) <= "00000011010000001100000000100110";
                        f_reg(123) <= "00100100001000100110000001100110";
                        f_reg(124) <= "00100101111100000110000001100110";
                        f_reg(125) <= "00010101001101110000000011001000";
                        f_reg(126) <= "10101100000010010000001100101100";
                        f_reg(127) <= "00110000001001001011001011011010";
                        f_reg(128) <= "00110001111100101011001011011010";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010101010110000000000011000010";
                        f_reg(132) <= "10101100000010100000001100110000";
                        f_reg(133) <= "00010101110111000000000011000000";
                        f_reg(134) <= "10101100000011100000001100110100";
                        f_reg(135) <= "00100100101001101010000010110001";
                        f_reg(136) <= "00100110011101001010000010110001";
                        f_reg(137) <= "00010100100100100000000010111100";
                        f_reg(138) <= "10101100000001000000001100111000";
                        f_reg(139) <= "00000000000000000000000000000000";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000110010000101100000000110";
                        f_reg(142) <= "00000010100101101100100000000110";
                        f_reg(143) <= "00111100000010011101000111110000";
                        f_reg(144) <= "00111100000101111101000111110000";
                        f_reg(145) <= "00010101011110010000000010110100";
                        f_reg(146) <= "10101100000010110000001100111100";
                        f_reg(147) <= "00101000011000011011011110100110";
                        f_reg(148) <= "00101010001011111011011110100110";
                        f_reg(149) <= "00101000101011101010010111101111";
                        f_reg(150) <= "00101010011111001010010111101111";
                        f_reg(151) <= "00010101110111000000000010101110";
                        f_reg(152) <= "10101100000011100000001101000000";
                        f_reg(153) <= "00111100000001000111001101000100";
                        f_reg(154) <= "00111100000100100111001101000100";
                        f_reg(155) <= "00000001010010010011000000100011";
                        f_reg(156) <= "00000011000101111010000000100011";
                        f_reg(157) <= "00000000000000000000000000000000";
                        f_reg(158) <= "00000000000000000000000000000000";
                        f_reg(159) <= "00000000010011000101100000000110";
                        f_reg(160) <= "00000010000110101100100000000110";
                        f_reg(161) <= "00010101000101100000000010100100";
                        f_reg(162) <= "10101100000010000000001101000100";
                        f_reg(163) <= "00000001011001110001100000100111";
                        f_reg(164) <= "00000011001101011000100000100111";
                        f_reg(165) <= "00010100111101010000000010100000";
                        f_reg(166) <= "10101100000001110000001101001000";
                        f_reg(167) <= "00010100011100010000000010011110";
                        f_reg(168) <= "10101100000000110000001101001100";
                        f_reg(169) <= "00000000100011010010100000101010";
                        f_reg(170) <= "00000010010110111001100000101010";
                        f_reg(171) <= "00000000110000010011000000100001";
                        f_reg(172) <= "00000010100011111010000000100001";
                        f_reg(173) <= "00010101000101100000000010011000";
                        f_reg(174) <= "10101100000010000000001101010000";
                        f_reg(175) <= "00000000000000000000000000000000";
                        f_reg(176) <= "00000000000000000000000000000000";
                        f_reg(177) <= "00000000000000000000000000000000";
                        f_reg(178) <= "00000000000000000000000000000000";
                        f_reg(179) <= "00000000000001010111000011000000";
                        f_reg(180) <= "00000000000100111110000011000000";
                        f_reg(181) <= "00000000000001010101001001000011";
                        f_reg(182) <= "00000000000100111100001001000011";
                        f_reg(183) <= "00100000110010011100101101101010";
                        f_reg(184) <= "00100010100101111100101101101010";
                        f_reg(185) <= "00010101110111000000000010001100";
                        f_reg(186) <= "10101100000011100000001101010100";
                        f_reg(187) <= "00010101010110000000000010001010";
                        f_reg(188) <= "10101100000010100000001101011000";
                        f_reg(189) <= "00010101001101110000000010001000";
                        f_reg(190) <= "10101100000010010000001101011100";
                        f_reg(191) <= "00010100110101000000000010000110";
                        f_reg(192) <= "10101100000001100000001101100000";
                        f_reg(193) <= "00100011110111011111111100000110";
                        f_reg(194) <= "00010011101000000000000000011000";
                        f_reg(195) <= "00100011110111011111111000001100";
                        f_reg(196) <= "00010011101000000000000000010110";
                        f_reg(197) <= "00100011110111011111110100010010";
                        f_reg(198) <= "00010011101000000000000000010100";
                        f_reg(199) <= "00100011110111101111111111111111";
                        f_reg(200) <= "00100011111111111111111111111111";
                        f_reg(201) <= "00010111110111110000000001111100";
                        f_reg(202) <= "00011111111000001111111101111101";
                        f_reg(203) <= "00010000000000000000000100000111";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000000000000000000000000000000";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00000000000000000000000000000000";
                        f_reg(215) <= "00000000000000000000000000000000";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "10001100000111010000011010111000";
                        f_reg(219) <= "00011111101000000000000000000011";
                        f_reg(220) <= "00100000000111010000000000111100";
                        f_reg(221) <= "00010000000000000000000000000010";
                        f_reg(222) <= "00100000000111010000000000000000";
                        f_reg(223) <= "00010100001011110000000001100110";
                        f_reg(224) <= "10101111101000010000011001000000";
                        f_reg(225) <= "10001100000111010000011010111000";
                        f_reg(226) <= "00011111101000000000000000000011";
                        f_reg(227) <= "00100000000111010000000000111100";
                        f_reg(228) <= "00010000000000000000000000000010";
                        f_reg(229) <= "00100000000111010000000000000000";
                        f_reg(230) <= "00010100010100000000000001011111";
                        f_reg(231) <= "10101111101000100000011001000100";
                        f_reg(232) <= "10001100000111010000011010111000";
                        f_reg(233) <= "00011111101000000000000000000011";
                        f_reg(234) <= "00100000000111010000000000111100";
                        f_reg(235) <= "00010000000000000000000000000010";
                        f_reg(236) <= "00100000000111010000000000000000";
                        f_reg(237) <= "00010100011100010000000001011000";
                        f_reg(238) <= "10101111101000110000011001001000";
                        f_reg(239) <= "10001100000111010000011010111000";
                        f_reg(240) <= "00011111101000000000000000000011";
                        f_reg(241) <= "00100000000111010000000000111100";
                        f_reg(242) <= "00010000000000000000000000000010";
                        f_reg(243) <= "00100000000111010000000000000000";
                        f_reg(244) <= "00010100100100100000000001010001";
                        f_reg(245) <= "10101111101001000000011001001100";
                        f_reg(246) <= "10001100000111010000011010111000";
                        f_reg(247) <= "00011111101000000000000000000011";
                        f_reg(248) <= "00100000000111010000000000111100";
                        f_reg(249) <= "00010000000000000000000000000010";
                        f_reg(250) <= "00100000000111010000000000000000";
                        f_reg(251) <= "00010100101100110000000001001010";
                        f_reg(252) <= "10101111101001010000011001010000";
                        f_reg(253) <= "10001100000111010000011010111000";
                        f_reg(254) <= "00011111101000000000000000000011";
                        f_reg(255) <= "00100000000111010000000000111100";
                        f_reg(256) <= "00010000000000000000000000000010";
                        f_reg(257) <= "00100000000111010000000000000000";
                        f_reg(258) <= "00010100110101000000000001000011";
                        f_reg(259) <= "10101111101001100000011001010100";
                        f_reg(260) <= "10001100000111010000011010111000";
                        f_reg(261) <= "00011111101000000000000000000011";
                        f_reg(262) <= "00100000000111010000000000111100";
                        f_reg(263) <= "00010000000000000000000000000010";
                        f_reg(264) <= "00100000000111010000000000000000";
                        f_reg(265) <= "00010100111101010000000000111100";
                        f_reg(266) <= "10101111101001110000011001011000";
                        f_reg(267) <= "10001100000111010000011010111000";
                        f_reg(268) <= "00011111101000000000000000000011";
                        f_reg(269) <= "00100000000111010000000000111100";
                        f_reg(270) <= "00010000000000000000000000000010";
                        f_reg(271) <= "00100000000111010000000000000000";
                        f_reg(272) <= "00010101000101100000000000110101";
                        f_reg(273) <= "10101111101010000000011001011100";
                        f_reg(274) <= "10001100000111010000011010111000";
                        f_reg(275) <= "00011111101000000000000000000011";
                        f_reg(276) <= "00100000000111010000000000111100";
                        f_reg(277) <= "00010000000000000000000000000010";
                        f_reg(278) <= "00100000000111010000000000000000";
                        f_reg(279) <= "00010101001101110000000000101110";
                        f_reg(280) <= "10101111101010010000011001100000";
                        f_reg(281) <= "10001100000111010000011010111000";
                        f_reg(282) <= "00011111101000000000000000000011";
                        f_reg(283) <= "00100000000111010000000000111100";
                        f_reg(284) <= "00010000000000000000000000000010";
                        f_reg(285) <= "00100000000111010000000000000000";
                        f_reg(286) <= "00010101010110000000000000100111";
                        f_reg(287) <= "10101111101010100000011001100100";
                        f_reg(288) <= "10001100000111010000011010111000";
                        f_reg(289) <= "00011111101000000000000000000011";
                        f_reg(290) <= "00100000000111010000000000111100";
                        f_reg(291) <= "00010000000000000000000000000010";
                        f_reg(292) <= "00100000000111010000000000000000";
                        f_reg(293) <= "00010101011110010000000000100000";
                        f_reg(294) <= "10101111101010110000011001101000";
                        f_reg(295) <= "10001100000111010000011010111000";
                        f_reg(296) <= "00011111101000000000000000000011";
                        f_reg(297) <= "00100000000111010000000000111100";
                        f_reg(298) <= "00010000000000000000000000000010";
                        f_reg(299) <= "00100000000111010000000000000000";
                        f_reg(300) <= "00010101100110100000000000011001";
                        f_reg(301) <= "10101111101011000000011001101100";
                        f_reg(302) <= "10001100000111010000011010111000";
                        f_reg(303) <= "00011111101000000000000000000011";
                        f_reg(304) <= "00100000000111010000000000111100";
                        f_reg(305) <= "00010000000000000000000000000010";
                        f_reg(306) <= "00100000000111010000000000000000";
                        f_reg(307) <= "00010101101110110000000000010010";
                        f_reg(308) <= "10101111101011010000011001110000";
                        f_reg(309) <= "10001100000111010000011010111000";
                        f_reg(310) <= "00011111101000000000000000000011";
                        f_reg(311) <= "00100000000111010000000000111100";
                        f_reg(312) <= "00010000000000000000000000000010";
                        f_reg(313) <= "00100000000111010000000000000000";
                        f_reg(314) <= "00010101110111000000000000001011";
                        f_reg(315) <= "10101111101011100000011001110100";
                        f_reg(316) <= "10001100000111010000011010111000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010111110111110000000000000100";
                        f_reg(322) <= "10101111101111100000011001111000";
                        f_reg(323) <= "10101100000111010000011010111000";
                        f_reg(324) <= "00010000000000001111111110000011";
                        f_reg(325) <= "10001100000111010000011010111000";
                        f_reg(326) <= "10001111101000010000011001000000";
                        f_reg(327) <= "10001100000111010000011010111000";
                        f_reg(328) <= "10001111101011110000011001000000";
                        f_reg(329) <= "00010100001011111111111111111100";
                        f_reg(330) <= "10001100000111010000011010111000";
                        f_reg(331) <= "10001111101000100000011001000100";
                        f_reg(332) <= "10001100000111010000011010111000";
                        f_reg(333) <= "10001111101100000000011001000100";
                        f_reg(334) <= "00010100010100001111111111111100";
                        f_reg(335) <= "10001100000111010000011010111000";
                        f_reg(336) <= "10001111101000110000011001001000";
                        f_reg(337) <= "10001100000111010000011010111000";
                        f_reg(338) <= "10001111101100010000011001001000";
                        f_reg(339) <= "00010100011100011111111111111100";
                        f_reg(340) <= "10001100000111010000011010111000";
                        f_reg(341) <= "10001111101001000000011001001100";
                        f_reg(342) <= "10001100000111010000011010111000";
                        f_reg(343) <= "10001111101100100000011001001100";
                        f_reg(344) <= "00010100100100101111111111111100";
                        f_reg(345) <= "10001100000111010000011010111000";
                        f_reg(346) <= "10001111101001010000011001010000";
                        f_reg(347) <= "10001100000111010000011010111000";
                        f_reg(348) <= "10001111101100110000011001010000";
                        f_reg(349) <= "00010100101100111111111111111100";
                        f_reg(350) <= "10001100000111010000011010111000";
                        f_reg(351) <= "10001111101001100000011001010100";
                        f_reg(352) <= "10001100000111010000011010111000";
                        f_reg(353) <= "10001111101101000000011001010100";
                        f_reg(354) <= "00010100110101001111111111111100";
                        f_reg(355) <= "10001100000111010000011010111000";
                        f_reg(356) <= "10001111101001110000011001011000";
                        f_reg(357) <= "10001100000111010000011010111000";
                        f_reg(358) <= "10001111101101010000011001011000";
                        f_reg(359) <= "00010100111101011111111111111100";
                        f_reg(360) <= "10001100000111010000011010111000";
                        f_reg(361) <= "10001111101010000000011001011100";
                        f_reg(362) <= "10001100000111010000011010111000";
                        f_reg(363) <= "10001111101101100000011001011100";
                        f_reg(364) <= "00010101000101101111111111111100";
                        f_reg(365) <= "10001100000111010000011010111000";
                        f_reg(366) <= "10001111101010010000011001100000";
                        f_reg(367) <= "10001100000111010000011010111000";
                        f_reg(368) <= "10001111101101110000011001100000";
                        f_reg(369) <= "00010101001101111111111111111100";
                        f_reg(370) <= "10001100000111010000011010111000";
                        f_reg(371) <= "10001111101010100000011001100100";
                        f_reg(372) <= "10001100000111010000011010111000";
                        f_reg(373) <= "10001111101110000000011001100100";
                        f_reg(374) <= "00010101010110001111111111111100";
                        f_reg(375) <= "10001100000111010000011010111000";
                        f_reg(376) <= "10001111101010110000011001101000";
                        f_reg(377) <= "10001100000111010000011010111000";
                        f_reg(378) <= "10001111101110010000011001101000";
                        f_reg(379) <= "00010101011110011111111111111100";
                        f_reg(380) <= "10001100000111010000011010111000";
                        f_reg(381) <= "10001111101011000000011001101100";
                        f_reg(382) <= "10001100000111010000011010111000";
                        f_reg(383) <= "10001111101110100000011001101100";
                        f_reg(384) <= "00010101100110101111111111111100";
                        f_reg(385) <= "10001100000111010000011010111000";
                        f_reg(386) <= "10001111101011010000011001110000";
                        f_reg(387) <= "10001100000111010000011010111000";
                        f_reg(388) <= "10001111101110110000011001110000";
                        f_reg(389) <= "00010101101110111111111111111100";
                        f_reg(390) <= "10001100000111010000011010111000";
                        f_reg(391) <= "10001111101011100000011001110100";
                        f_reg(392) <= "10001100000111010000011010111000";
                        f_reg(393) <= "10001111101111000000011001110100";
                        f_reg(394) <= "00010101110111001111111111111100";
                        f_reg(395) <= "10001100000111010000011010111000";
                        f_reg(396) <= "10001111101111100000011001111000";
                        f_reg(397) <= "10001100000111010000011010111000";
                        f_reg(398) <= "10001111101111110000011001111000";
                        f_reg(399) <= "00010111110111111111111111111100";
                        f_reg(400) <= "00010000000000001111111100110111";
                        f_reg(401) <= "00000000000000000000000000000000";
                        f_reg(402) <= "00000000000000000000000000000000";
                        f_reg(403) <= "00000000000000000000000000000000";
                        f_reg(404) <= "00000000000000000000000000000000";
                        f_reg(405) <= "00000000000000000000000000000000";
                        f_reg(406) <= "00000000000000000000000000000000";
                        f_reg(407) <= "00000000000000000000000000000000";
                        f_reg(408) <= "00000000000000000000000000000000";
                        f_reg(409) <= "00000000000000000000000000000000";
                        f_reg(410) <= "00000000000000000000000000000000";
                        f_reg(411) <= "00000000000000000000000000000000";
                        f_reg(412) <= "00000000000000000000000000000000";
                        f_reg(413) <= "00000000000000000000000000000000";
                        f_reg(414) <= "00000000000000000000000000000000";
                        f_reg(415) <= "00000000000000000000000000000000";
                        f_reg(416) <= "00000000000000000000000000000000";
                        f_reg(417) <= "00000000000000000000000000000000";
                        f_reg(418) <= "00000000000000000000000000000000";
                        f_reg(419) <= "00000000000000000000000000000000";
                        f_reg(420) <= "00000000000000000000000000000000";
                        f_reg(421) <= "00000000000000000000000000000000";
                        f_reg(422) <= "00000000000000000000000000000000";
                        f_reg(423) <= "00000000000000000000000000000000";
                        f_reg(424) <= "00000000000000000000000000000000";
                        f_reg(425) <= "00000000000000000000000000000000";
                        f_reg(426) <= "00000000000000000000000000000000";
                        f_reg(427) <= "00000000000000000000000000000000";
                        f_reg(428) <= "00000000000000000000000000000000";
                        f_reg(429) <= "00000000000000000000000000000000";
                        f_reg(430) <= "00000000000000000000000000000000";
                        f_reg(431) <= "00000000000000000000001111100111";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 -31521
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SLTI R2 R0 5593
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SLTIU R3 R0 2299
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SLLV R4 R0 R2
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SUBU R5 R2 R0
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- ADD R6 R2 R5
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- SLT R7 R4 R4
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- ADDU R8 R7 R4
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- SLTIU R9 R0 -17025
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- NOR R10 R8 R0
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- AND R11 R10 R9
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- ADDIU R12 R7 27880
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- ADDI R13 R5 32229
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- SLTI R14 R6 4484
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- ORI R15 R5 21919
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- OR R16 R8 R8
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SUB R17 R8 R0
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- ADDU R18 R15 R13
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SLLV R19 R1 R7
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- ADD R20 R5 R14
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- ADD R21 R16 R19
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- NOP
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- ADDI R22 R4 -29515
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- NOP
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- SUB R23 R18 R11
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- XOR R24 R12 R0
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- ADDIU R25 R20 24678
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- SW R17 R0 812
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- ANDI R26 R20 -19750
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- NOP
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- SW R24 R0 816
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- SW R23 R0 820
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- ADDIU R27 R22 -24399
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- SW R26 R0 824
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- NOP
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- SRLV R28 R8 R27
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- LUI R29 -11792
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- SW R28 R0 828
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- SLTI R30 R3 -18522
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- SLTI R2 R22 -23057
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SW R2 R0 832
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- LUI R10 29508
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- SUBU R9 R24 R29
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- NOP
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- SRLV R6 R12 R25
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- SW R8 R0 836
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- NOR R15 R6 R21
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- SW R21 R0 840
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SW R15 R0 844
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- SLT R1 R10 R13
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- ADDU R9 R9 R30
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SW R8 R0 848
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- NOP
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- NOP
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SLL R7 R1 3
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- SRA R5 R1 9
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- ADDI R14 R9 -13462
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SW R7 R0 852
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- SW R5 R0 856
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- SW R14 R0 860
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- SW R9 R0 864
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- ADDI R31 R31 -1
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- BGTZ R31 -62
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- BEQ R0 R0 400
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- LUI R30 999
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- LUI R31 999
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- SRL R30 R30 16
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SRL R31 R31 16
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- LUI R1 -31521
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- LUI R15 -31521
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SLTI R2 R0 5593
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- SLTI R16 R0 5593
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- SLTIU R3 R0 2299
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- SLTIU R17 R0 2299
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- SLLV R4 R0 R2
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- SLLV R18 R0 R16
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- SUBU R5 R2 R0
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- SUBU R19 R16 R0
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- ADD R6 R2 R5
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- ADD R20 R16 R19
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SLT R7 R4 R4
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- SLT R21 R18 R18
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- ADDU R8 R7 R4
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- ADDU R22 R21 R18
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SLTIU R9 R0 -17025
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- SLTIU R23 R0 -17025
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- NOR R10 R8 R0
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- NOR R24 R22 R0
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- AND R11 R10 R9
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- AND R25 R24 R23
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- ADDIU R12 R7 27880
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- ADDIU R26 R21 27880
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- ADDI R13 R5 32229
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- ADDI R27 R19 32229
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SLTI R14 R6 4484
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SLTI R28 R20 4484
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- ORI R2 R5 21919
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- ORI R16 R19 21919
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- OR R10 R8 R8
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- OR R24 R22 R22
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SUB R9 R8 R0
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- SUB R23 R22 R0
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- ADDU R6 R2 R13
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- ADDU R20 R16 R27
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- SLLV R2 R1 R7
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- SLLV R16 R15 R21
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- ADD R1 R5 R14
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- ADD R15 R19 R28
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- ADD R7 R10 R2
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- ADD R21 R24 R16
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- NOP
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- NOP
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- ADDI R5 R4 -29515
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- ADDI R19 R18 -29515
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- NOP
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- NOP
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- SUB R14 R6 R11
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- SUB R28 R20 R25
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- XOR R10 R12 R0
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- XOR R24 R26 R0
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- ADDIU R2 R1 24678
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- ADDIU R16 R15 24678
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- BNE R9 R23 200
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- SW R9 R0 812
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- ANDI R4 R1 -19750
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- ANDI R18 R15 -19750
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- NOP
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- NOP
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- BNE R10 R24 194
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- SW R10 R0 816
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- BNE R14 R28 192
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- SW R14 R0 820
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- ADDIU R6 R5 -24399
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- ADDIU R20 R19 -24399
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- BNE R4 R18 188
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SW R4 R0 824
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- NOP
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- NOP
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- SRLV R11 R8 R6
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- SRLV R25 R22 R20
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- LUI R9 -11792
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- LUI R23 -11792
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- BNE R11 R25 180
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- SW R11 R0 828
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- SLTI R1 R3 -18522
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- SLTI R15 R17 -18522
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- SLTI R14 R5 -23057
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- SLTI R28 R19 -23057
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- BNE R14 R28 174
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- SW R14 R0 832
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- LUI R4 29508
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- LUI R18 29508
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- SUBU R6 R10 R9
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- SUBU R20 R24 R23
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- NOP
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- NOP
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- SRLV R11 R12 R2
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- SRLV R25 R26 R16
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- BNE R8 R22 164
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- SW R8 R0 836
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- NOR R3 R11 R7
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- NOR R17 R25 R21
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- BNE R7 R21 160
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- SW R7 R0 840
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- BNE R3 R17 158
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- SW R3 R0 844
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- SLT R5 R4 R13
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- SLT R19 R18 R27
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- ADDU R6 R6 R1
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- ADDU R20 R20 R15
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- BNE R8 R22 152
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- SW R8 R0 848
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- NOP
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- NOP
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- NOP
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- NOP
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- SLL R14 R5 3
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- SLL R28 R19 3
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- SRA R10 R5 9
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SRA R24 R19 9
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- ADDI R9 R6 -13462
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- ADDI R23 R20 -13462
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- BNE R14 R28 140
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- SW R14 R0 852
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- BNE R10 R24 138
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- SW R10 R0 856
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- BNE R9 R23 136
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- SW R9 R0 860
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- BNE R6 R20 134
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- SW R6 R0 864
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- ADDI R29 R30 -250
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- BEQ R29 R0 24
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- ADDI R29 R30 -500
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- BEQ R29 R0 22
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- ADDI R29 R30 -750
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- BEQ R29 R0 20
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- ADDI R30 R30 -1
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- ADDI R31 R31 -1
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- BNE R30 R31 124
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- BGTZ R31 -131
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- BEQ R0 R0 263
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- NOP
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- NOP
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- NOP
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- NOP
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- NOP
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- NOP
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- NOP
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- NOP
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- NOP
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- NOP
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- NOP
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- NOP
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- NOP
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- NOP
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- LW R29 R0 1720
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- BGTZ R29 3
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- ADDI R29 R0 60
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- BEQ R0 R0 2
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- ADDI R29 R0 0
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- BNE R1 R15 102
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- SW R1 R29 1600
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- LW R29 R0 1720
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- BGTZ R29 3
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- ADDI R29 R0 60
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- BEQ R0 R0 2
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- ADDI R29 R0 0
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- BNE R2 R16 95
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- SW R2 R29 1604
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- LW R29 R0 1720
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- BGTZ R29 3
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- ADDI R29 R0 60
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- BEQ R0 R0 2
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- ADDI R29 R0 0
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- BNE R3 R17 88
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- SW R3 R29 1608
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- LW R29 R0 1720
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- BGTZ R29 3
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- ADDI R29 R0 60
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- BEQ R0 R0 2
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- ADDI R29 R0 0
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- BNE R4 R18 81
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- SW R4 R29 1612
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- LW R29 R0 1720
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- BGTZ R29 3
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- ADDI R29 R0 60
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- BEQ R0 R0 2
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- ADDI R29 R0 0
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- BNE R5 R19 74
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- SW R5 R29 1616
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- LW R29 R0 1720
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- BGTZ R29 3
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- ADDI R29 R0 60
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- BEQ R0 R0 2
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- ADDI R29 R0 0
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- BNE R6 R20 67
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- SW R6 R29 1620
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- LW R29 R0 1720
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- BGTZ R29 3
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- ADDI R29 R0 60
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- BEQ R0 R0 2
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- ADDI R29 R0 0
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- BNE R7 R21 60
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- SW R7 R29 1624
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- LW R29 R0 1720
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- BGTZ R29 3
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- ADDI R29 R0 60
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- BEQ R0 R0 2
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- ADDI R29 R0 0
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- BNE R8 R22 53
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- SW R8 R29 1628
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- LW R29 R0 1720
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- BGTZ R29 3
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- ADDI R29 R0 60
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- BEQ R0 R0 2
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- ADDI R29 R0 0
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- BNE R9 R23 46
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- SW R9 R29 1632
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- LW R29 R0 1720
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- BGTZ R29 3
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- ADDI R29 R0 60
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- BEQ R0 R0 2
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- ADDI R29 R0 0
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- BNE R10 R24 39
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- SW R10 R29 1636
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- LW R29 R0 1720
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- BGTZ R29 3
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- ADDI R29 R0 60
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- BEQ R0 R0 2
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- ADDI R29 R0 0
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- BNE R11 R25 32
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- SW R11 R29 1640
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- LW R29 R0 1720
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- BGTZ R29 3
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- ADDI R29 R0 60
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- BEQ R0 R0 2
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- ADDI R29 R0 0
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- BNE R12 R26 25
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- SW R12 R29 1644
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- LW R29 R0 1720
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- BGTZ R29 3
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- ADDI R29 R0 60
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- BEQ R0 R0 2
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- ADDI R29 R0 0
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- BNE R13 R27 18
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- SW R13 R29 1648
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- LW R29 R0 1720
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- BGTZ R29 3
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- ADDI R29 R0 60
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- BEQ R0 R0 2
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- ADDI R29 R0 0
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- BNE R14 R28 11
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- SW R14 R29 1652
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- LW R29 R0 1720
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- BGTZ R29 3
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- ADDI R29 R0 60
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- BEQ R0 R0 2
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- ADDI R29 R0 0
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- BNE R30 R31 4
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- SW R30 R29 1656
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- SW R29 R0 1720
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- BEQ R0 R0 -125
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- LW R29 R0 1720
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- LW R1 R29 1600
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- LW R29 R0 1720
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- LW R15 R29 1600
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- BNE R1 R15 -4
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- LW R29 R0 1720
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- LW R2 R29 1604
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- LW R29 R0 1720
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- LW R16 R29 1604
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- BNE R2 R16 -4
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- LW R29 R0 1720
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- LW R3 R29 1608
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- LW R29 R0 1720
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- LW R17 R29 1608
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- BNE R3 R17 -4
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- LW R29 R0 1720
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- LW R4 R29 1612
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- LW R29 R0 1720
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- LW R18 R29 1612
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- BNE R4 R18 -4
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- LW R29 R0 1720
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- LW R5 R29 1616
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- LW R29 R0 1720
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- LW R19 R29 1616
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- BNE R5 R19 -4
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- LW R29 R0 1720
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- LW R6 R29 1620
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- LW R29 R0 1720
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- LW R20 R29 1620
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- BNE R6 R20 -4
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- LW R29 R0 1720
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- LW R7 R29 1624
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- LW R29 R0 1720
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- LW R21 R29 1624
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- BNE R7 R21 -4
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- LW R29 R0 1720
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- LW R8 R29 1628
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- LW R29 R0 1720
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- LW R22 R29 1628
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- BNE R8 R22 -4
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- LW R29 R0 1720
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- LW R9 R29 1632
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- LW R29 R0 1720
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- LW R23 R29 1632
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- BNE R9 R23 -4
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- LW R29 R0 1720
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- LW R10 R29 1636
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- LW R29 R0 1720
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- LW R24 R29 1636
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- BNE R10 R24 -4
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- LW R29 R0 1720
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- LW R11 R29 1640
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- LW R29 R0 1720
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- LW R25 R29 1640
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- BNE R11 R25 -4
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- LW R29 R0 1720
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- LW R12 R29 1644
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- LW R29 R0 1720
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- LW R26 R29 1644
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- BNE R12 R26 -4
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- LW R29 R0 1720
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- LW R13 R29 1648
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- LW R29 R0 1720
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- LW R27 R29 1648
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- BNE R13 R27 -4
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- LW R29 R0 1720
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- LW R14 R29 1652
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- LW R29 R0 1720
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- LW R28 R29 1652
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- BNE R14 R28 -4
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- LW R29 R0 1720
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- LW R30 R29 1656
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- LW R29 R0 1720
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- LW R31 R29 1656
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- BNE R30 R31 -4
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- BEQ R0 R0 -201
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- NOP
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- NOP
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- NOP
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- NOP
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- NOP
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- NOP
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- NOP
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- NOP
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- NOP
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- NOP
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- NOP
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- NOP
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- NOP
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- NOP
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- NOP
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- NOP
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- NOP
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- NOP
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- NOP
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- NOP
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- NOP
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- NOP
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- NOP
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- NOP
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- NOP
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- NOP
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- NOP
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- NOP
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- NOP
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- NOP
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- NOP
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- NOP
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- NOP
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- NOP
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- NOP
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- NOP
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- NOP
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- NOP
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- NOP
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- NOP
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- NOP
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- NOP
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- NOP
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- NOP
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- NOP
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- NOP
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- NOP
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- NOP
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- NOP
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- NOP
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- NOP
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- NOP
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- NOP
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- NOP
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- NOP
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- NOP
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- NOP
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- NOP
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- NOP
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- NOP
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- NOP
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- NOP
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- NOP
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- NOP
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- NOP
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011000010011011111";
                        f_reg(4) <= "00101000000000100001010111011001";
                        f_reg(5) <= "00101100000000110000100011111011";
                        f_reg(6) <= "00000000010000000010000000000100";
                        f_reg(7) <= "00000000010000000010100000100011";
                        f_reg(8) <= "00000000010001010011000000100000";
                        f_reg(9) <= "00000000100001000011100000101010";
                        f_reg(10) <= "00000000111001000100000000100001";
                        f_reg(11) <= "00101100000010011011110101111111";
                        f_reg(12) <= "00000001000000000101000000100111";
                        f_reg(13) <= "00000001010010010101100000100100";
                        f_reg(14) <= "00100100111011000110110011101000";
                        f_reg(15) <= "00100000101011010111110111100101";
                        f_reg(16) <= "00101000110011100001000110000100";
                        f_reg(17) <= "00110100101011110101010110011111";
                        f_reg(18) <= "00000001000010001000000000100101";
                        f_reg(19) <= "00000001000000001000100000100010";
                        f_reg(20) <= "00000001111011011001000000100001";
                        f_reg(21) <= "00000000111000011001100000000100";
                        f_reg(22) <= "00000000101011101010000000100000";
                        f_reg(23) <= "00000010000100111010100000100000";
                        f_reg(24) <= "00000000000000000000000000000000";
                        f_reg(25) <= "00100000100101101000110010110101";
                        f_reg(26) <= "00000000000000000000000000000000";
                        f_reg(27) <= "00000010010010111011100000100010";
                        f_reg(28) <= "00000001100000001100000000100110";
                        f_reg(29) <= "00100110100110010110000001100110";
                        f_reg(30) <= "10101100000100010000001100101100";
                        f_reg(31) <= "00110010100110101011001011011010";
                        f_reg(32) <= "00000000000000000000000000000000";
                        f_reg(33) <= "10101100000110000000001100110000";
                        f_reg(34) <= "10101100000101110000001100110100";
                        f_reg(35) <= "00100110110110111010000010110001";
                        f_reg(36) <= "10101100000110100000001100111000";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00000011011010001110000000000110";
                        f_reg(39) <= "00111100000111011101000111110000";
                        f_reg(40) <= "10101100000111000000001100111100";
                        f_reg(41) <= "00101000011111101011011110100110";
                        f_reg(42) <= "00101010110000101010010111101111";
                        f_reg(43) <= "10101100000000100000001101000000";
                        f_reg(44) <= "00111100000010100111001101000100";
                        f_reg(45) <= "00000011000111010100100000100011";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00000011001011000011000000000110";
                        f_reg(48) <= "10101100000010000000001101000100";
                        f_reg(49) <= "00000000110101010111100000100111";
                        f_reg(50) <= "10101100000101010000001101001000";
                        f_reg(51) <= "10101100000011110000001101001100";
                        f_reg(52) <= "00000001010011010000100000101010";
                        f_reg(53) <= "00000001001111100100100000100001";
                        f_reg(54) <= "10101100000010000000001101010000";
                        f_reg(55) <= "00000000000000000000000000000000";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000010011100011000000";
                        f_reg(58) <= "00000000000000010010101001000011";
                        f_reg(59) <= "00100001001011101100101101101010";
                        f_reg(60) <= "10101100000001110000001101010100";
                        f_reg(61) <= "10101100000001010000001101011000";
                        f_reg(62) <= "10101100000011100000001101011100";
                        f_reg(63) <= "10101100000010010000001101100000";
                        f_reg(64) <= "00100011111111111111111111111111";
                        f_reg(65) <= "00011111111000001111111111000010";
                        f_reg(66) <= "00010000000000000000000110010000";
                        f_reg(67) <= "00111100000111100000001111100111";
                        f_reg(68) <= "00111100000111110000001111100111";
                        f_reg(69) <= "00000000000111101111010000000010";
                        f_reg(70) <= "00000000000111111111110000000010";
                        f_reg(71) <= "00111100000000011000010011011111";
                        f_reg(72) <= "00111100000011111000010011011111";
                        f_reg(73) <= "00101000000000100001010111011001";
                        f_reg(74) <= "00101000000100000001010111011001";
                        f_reg(75) <= "00101100000000110000100011111011";
                        f_reg(76) <= "00101100000100010000100011111011";
                        f_reg(77) <= "00000000010000000010000000000100";
                        f_reg(78) <= "00000010000000001001000000000100";
                        f_reg(79) <= "00000000010000000010100000100011";
                        f_reg(80) <= "00000010000000001001100000100011";
                        f_reg(81) <= "00000000010001010011000000100000";
                        f_reg(82) <= "00000010000100111010000000100000";
                        f_reg(83) <= "00000000100001000011100000101010";
                        f_reg(84) <= "00000010010100101010100000101010";
                        f_reg(85) <= "00000000111001000100000000100001";
                        f_reg(86) <= "00000010101100101011000000100001";
                        f_reg(87) <= "00101100000010011011110101111111";
                        f_reg(88) <= "00101100000101111011110101111111";
                        f_reg(89) <= "00000001000000000101000000100111";
                        f_reg(90) <= "00000010110000001100000000100111";
                        f_reg(91) <= "00000001010010010101100000100100";
                        f_reg(92) <= "00000011000101111100100000100100";
                        f_reg(93) <= "00100100111011000110110011101000";
                        f_reg(94) <= "00100110101110100110110011101000";
                        f_reg(95) <= "00100000101011010111110111100101";
                        f_reg(96) <= "00100010011110110111110111100101";
                        f_reg(97) <= "00101000110011100001000110000100";
                        f_reg(98) <= "00101010100111000001000110000100";
                        f_reg(99) <= "00110100101000100101010110011111";
                        f_reg(100) <= "00110110011100000101010110011111";
                        f_reg(101) <= "00000001000010000101000000100101";
                        f_reg(102) <= "00000010110101101100000000100101";
                        f_reg(103) <= "00000001000000000100100000100010";
                        f_reg(104) <= "00000010110000001011100000100010";
                        f_reg(105) <= "00000000010011010011000000100001";
                        f_reg(106) <= "00000010000110111010000000100001";
                        f_reg(107) <= "00000000111000010001000000000100";
                        f_reg(108) <= "00000010101011111000000000000100";
                        f_reg(109) <= "00000000101011100000100000100000";
                        f_reg(110) <= "00000010011111000111100000100000";
                        f_reg(111) <= "00000001010000100011100000100000";
                        f_reg(112) <= "00000011000100001010100000100000";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00100000100001011000110010110101";
                        f_reg(116) <= "00100010010100111000110010110101";
                        f_reg(117) <= "00000000000000000000000000000000";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000110010110111000000100010";
                        f_reg(120) <= "00000010100110011110000000100010";
                        f_reg(121) <= "00000001100000000101000000100110";
                        f_reg(122) <= "00000011010000001100000000100110";
                        f_reg(123) <= "00100100001000100110000001100110";
                        f_reg(124) <= "00100101111100000110000001100110";
                        f_reg(125) <= "00010101001101110000000011001000";
                        f_reg(126) <= "10101100000010010000001100101100";
                        f_reg(127) <= "00110000001001001011001011011010";
                        f_reg(128) <= "00110001111100101011001011011010";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010101010110000000000011000010";
                        f_reg(132) <= "10101100000010100000001100110000";
                        f_reg(133) <= "00010101110111000000000011000000";
                        f_reg(134) <= "10101100000011100000001100110100";
                        f_reg(135) <= "00100100101001101010000010110001";
                        f_reg(136) <= "00100110011101001010000010110001";
                        f_reg(137) <= "00010100100100100000000010111100";
                        f_reg(138) <= "10101100000001000000001100111000";
                        f_reg(139) <= "00000000000000000000000000000000";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000110010000101100000000110";
                        f_reg(142) <= "00000010100101101100100000000110";
                        f_reg(143) <= "00111100000010011101000111110000";
                        f_reg(144) <= "00111100000101111101000111110000";
                        f_reg(145) <= "00010101011110010000000010110100";
                        f_reg(146) <= "10101100000010110000001100111100";
                        f_reg(147) <= "00101000011000011011011110100110";
                        f_reg(148) <= "00101010001011111011011110100110";
                        f_reg(149) <= "00101000101011101010010111101111";
                        f_reg(150) <= "00101010011111001010010111101111";
                        f_reg(151) <= "00010101110111000000000010101110";
                        f_reg(152) <= "10101100000011100000001101000000";
                        f_reg(153) <= "00111100000001000111001101000100";
                        f_reg(154) <= "00111100000100100111001101000100";
                        f_reg(155) <= "00000001010010010011000000100011";
                        f_reg(156) <= "00000011000101111010000000100011";
                        f_reg(157) <= "00000000000000000000000000000000";
                        f_reg(158) <= "00000000000000000000000000000000";
                        f_reg(159) <= "00000000010011000101100000000110";
                        f_reg(160) <= "00000010000110101100100000000110";
                        f_reg(161) <= "00010101000101100000000010100100";
                        f_reg(162) <= "10101100000010000000001101000100";
                        f_reg(163) <= "00000001011001110001100000100111";
                        f_reg(164) <= "00000011001101011000100000100111";
                        f_reg(165) <= "00010100111101010000000010100000";
                        f_reg(166) <= "10101100000001110000001101001000";
                        f_reg(167) <= "00010100011100010000000010011110";
                        f_reg(168) <= "10101100000000110000001101001100";
                        f_reg(169) <= "00000000100011010010100000101010";
                        f_reg(170) <= "00000010010110111001100000101010";
                        f_reg(171) <= "00000000110000010011000000100001";
                        f_reg(172) <= "00000010100011111010000000100001";
                        f_reg(173) <= "00010101000101100000000010011000";
                        f_reg(174) <= "10101100000010000000001101010000";
                        f_reg(175) <= "00000000000000000000000000000000";
                        f_reg(176) <= "00000000000000000000000000000000";
                        f_reg(177) <= "00000000000000000000000000000000";
                        f_reg(178) <= "00000000000000000000000000000000";
                        f_reg(179) <= "00000000000001010111000011000000";
                        f_reg(180) <= "00000000000100111110000011000000";
                        f_reg(181) <= "00000000000001010101001001000011";
                        f_reg(182) <= "00000000000100111100001001000011";
                        f_reg(183) <= "00100000110010011100101101101010";
                        f_reg(184) <= "00100010100101111100101101101010";
                        f_reg(185) <= "00010101110111000000000010001100";
                        f_reg(186) <= "10101100000011100000001101010100";
                        f_reg(187) <= "00010101010110000000000010001010";
                        f_reg(188) <= "10101100000010100000001101011000";
                        f_reg(189) <= "00010101001101110000000010001000";
                        f_reg(190) <= "10101100000010010000001101011100";
                        f_reg(191) <= "00010100110101000000000010000110";
                        f_reg(192) <= "10101100000001100000001101100000";
                        f_reg(193) <= "00100011110111011111111100000110";
                        f_reg(194) <= "00010011101000000000000000011000";
                        f_reg(195) <= "00100011110111011111111000001100";
                        f_reg(196) <= "00010011101000000000000000010110";
                        f_reg(197) <= "00100011110111011111110100010010";
                        f_reg(198) <= "00010011101000000000000000010100";
                        f_reg(199) <= "00100011110111101111111111111111";
                        f_reg(200) <= "00100011111111111111111111111111";
                        f_reg(201) <= "00010111110111110000000001111100";
                        f_reg(202) <= "00011111111000001111111101111101";
                        f_reg(203) <= "00010000000000000000000100000111";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000000000000000000000000000000";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00000000000000000000000000000000";
                        f_reg(215) <= "00000000000000000000000000000000";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "10001100000111010000011010111000";
                        f_reg(219) <= "00011111101000000000000000000011";
                        f_reg(220) <= "00100000000111010000000000111100";
                        f_reg(221) <= "00010000000000000000000000000010";
                        f_reg(222) <= "00100000000111010000000000000000";
                        f_reg(223) <= "00010100001011110000000001100110";
                        f_reg(224) <= "10101111101000010000011001000000";
                        f_reg(225) <= "10001100000111010000011010111000";
                        f_reg(226) <= "00011111101000000000000000000011";
                        f_reg(227) <= "00100000000111010000000000111100";
                        f_reg(228) <= "00010000000000000000000000000010";
                        f_reg(229) <= "00100000000111010000000000000000";
                        f_reg(230) <= "00010100010100000000000001011111";
                        f_reg(231) <= "10101111101000100000011001000100";
                        f_reg(232) <= "10001100000111010000011010111000";
                        f_reg(233) <= "00011111101000000000000000000011";
                        f_reg(234) <= "00100000000111010000000000111100";
                        f_reg(235) <= "00010000000000000000000000000010";
                        f_reg(236) <= "00100000000111010000000000000000";
                        f_reg(237) <= "00010100011100010000000001011000";
                        f_reg(238) <= "10101111101000110000011001001000";
                        f_reg(239) <= "10001100000111010000011010111000";
                        f_reg(240) <= "00011111101000000000000000000011";
                        f_reg(241) <= "00100000000111010000000000111100";
                        f_reg(242) <= "00010000000000000000000000000010";
                        f_reg(243) <= "00100000000111010000000000000000";
                        f_reg(244) <= "00010100100100100000000001010001";
                        f_reg(245) <= "10101111101001000000011001001100";
                        f_reg(246) <= "10001100000111010000011010111000";
                        f_reg(247) <= "00011111101000000000000000000011";
                        f_reg(248) <= "00100000000111010000000000111100";
                        f_reg(249) <= "00010000000000000000000000000010";
                        f_reg(250) <= "00100000000111010000000000000000";
                        f_reg(251) <= "00010100101100110000000001001010";
                        f_reg(252) <= "10101111101001010000011001010000";
                        f_reg(253) <= "10001100000111010000011010111000";
                        f_reg(254) <= "00011111101000000000000000000011";
                        f_reg(255) <= "00100000000111010000000000111100";
                        f_reg(256) <= "00010000000000000000000000000010";
                        f_reg(257) <= "00100000000111010000000000000000";
                        f_reg(258) <= "00010100110101000000000001000011";
                        f_reg(259) <= "10101111101001100000011001010100";
                        f_reg(260) <= "10001100000111010000011010111000";
                        f_reg(261) <= "00011111101000000000000000000011";
                        f_reg(262) <= "00100000000111010000000000111100";
                        f_reg(263) <= "00010000000000000000000000000010";
                        f_reg(264) <= "00100000000111010000000000000000";
                        f_reg(265) <= "00010100111101010000000000111100";
                        f_reg(266) <= "10101111101001110000011001011000";
                        f_reg(267) <= "10001100000111010000011010111000";
                        f_reg(268) <= "00011111101000000000000000000011";
                        f_reg(269) <= "00100000000111010000000000111100";
                        f_reg(270) <= "00010000000000000000000000000010";
                        f_reg(271) <= "00100000000111010000000000000000";
                        f_reg(272) <= "00010101000101100000000000110101";
                        f_reg(273) <= "10101111101010000000011001011100";
                        f_reg(274) <= "10001100000111010000011010111000";
                        f_reg(275) <= "00011111101000000000000000000011";
                        f_reg(276) <= "00100000000111010000000000111100";
                        f_reg(277) <= "00010000000000000000000000000010";
                        f_reg(278) <= "00100000000111010000000000000000";
                        f_reg(279) <= "00010101001101110000000000101110";
                        f_reg(280) <= "10101111101010010000011001100000";
                        f_reg(281) <= "10001100000111010000011010111000";
                        f_reg(282) <= "00011111101000000000000000000011";
                        f_reg(283) <= "00100000000111010000000000111100";
                        f_reg(284) <= "00010000000000000000000000000010";
                        f_reg(285) <= "00100000000111010000000000000000";
                        f_reg(286) <= "00010101010110000000000000100111";
                        f_reg(287) <= "10101111101010100000011001100100";
                        f_reg(288) <= "10001100000111010000011010111000";
                        f_reg(289) <= "00011111101000000000000000000011";
                        f_reg(290) <= "00100000000111010000000000111100";
                        f_reg(291) <= "00010000000000000000000000000010";
                        f_reg(292) <= "00100000000111010000000000000000";
                        f_reg(293) <= "00010101011110010000000000100000";
                        f_reg(294) <= "10101111101010110000011001101000";
                        f_reg(295) <= "10001100000111010000011010111000";
                        f_reg(296) <= "00011111101000000000000000000011";
                        f_reg(297) <= "00100000000111010000000000111100";
                        f_reg(298) <= "00010000000000000000000000000010";
                        f_reg(299) <= "00100000000111010000000000000000";
                        f_reg(300) <= "00010101100110100000000000011001";
                        f_reg(301) <= "10101111101011000000011001101100";
                        f_reg(302) <= "10001100000111010000011010111000";
                        f_reg(303) <= "00011111101000000000000000000011";
                        f_reg(304) <= "00100000000111010000000000111100";
                        f_reg(305) <= "00010000000000000000000000000010";
                        f_reg(306) <= "00100000000111010000000000000000";
                        f_reg(307) <= "00010101101110110000000000010010";
                        f_reg(308) <= "10101111101011010000011001110000";
                        f_reg(309) <= "10001100000111010000011010111000";
                        f_reg(310) <= "00011111101000000000000000000011";
                        f_reg(311) <= "00100000000111010000000000111100";
                        f_reg(312) <= "00010000000000000000000000000010";
                        f_reg(313) <= "00100000000111010000000000000000";
                        f_reg(314) <= "00010101110111000000000000001011";
                        f_reg(315) <= "10101111101011100000011001110100";
                        f_reg(316) <= "10001100000111010000011010111000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010111110111110000000000000100";
                        f_reg(322) <= "10101111101111100000011001111000";
                        f_reg(323) <= "10101100000111010000011010111000";
                        f_reg(324) <= "00010000000000001111111110000011";
                        f_reg(325) <= "10001100000111010000011010111000";
                        f_reg(326) <= "10001111101000010000011001000000";
                        f_reg(327) <= "10001100000111010000011010111000";
                        f_reg(328) <= "10001111101011110000011001000000";
                        f_reg(329) <= "00010100001011111111111111111100";
                        f_reg(330) <= "10001100000111010000011010111000";
                        f_reg(331) <= "10001111101000100000011001000100";
                        f_reg(332) <= "10001100000111010000011010111000";
                        f_reg(333) <= "10001111101100000000011001000100";
                        f_reg(334) <= "00010100010100001111111111111100";
                        f_reg(335) <= "10001100000111010000011010111000";
                        f_reg(336) <= "10001111101000110000011001001000";
                        f_reg(337) <= "10001100000111010000011010111000";
                        f_reg(338) <= "10001111101100010000011001001000";
                        f_reg(339) <= "00010100011100011111111111111100";
                        f_reg(340) <= "10001100000111010000011010111000";
                        f_reg(341) <= "10001111101001000000011001001100";
                        f_reg(342) <= "10001100000111010000011010111000";
                        f_reg(343) <= "10001111101100100000011001001100";
                        f_reg(344) <= "00010100100100101111111111111100";
                        f_reg(345) <= "10001100000111010000011010111000";
                        f_reg(346) <= "10001111101001010000011001010000";
                        f_reg(347) <= "10001100000111010000011010111000";
                        f_reg(348) <= "10001111101100110000011001010000";
                        f_reg(349) <= "00010100101100111111111111111100";
                        f_reg(350) <= "10001100000111010000011010111000";
                        f_reg(351) <= "10001111101001100000011001010100";
                        f_reg(352) <= "10001100000111010000011010111000";
                        f_reg(353) <= "10001111101101000000011001010100";
                        f_reg(354) <= "00010100110101001111111111111100";
                        f_reg(355) <= "10001100000111010000011010111000";
                        f_reg(356) <= "10001111101001110000011001011000";
                        f_reg(357) <= "10001100000111010000011010111000";
                        f_reg(358) <= "10001111101101010000011001011000";
                        f_reg(359) <= "00010100111101011111111111111100";
                        f_reg(360) <= "10001100000111010000011010111000";
                        f_reg(361) <= "10001111101010000000011001011100";
                        f_reg(362) <= "10001100000111010000011010111000";
                        f_reg(363) <= "10001111101101100000011001011100";
                        f_reg(364) <= "00010101000101101111111111111100";
                        f_reg(365) <= "10001100000111010000011010111000";
                        f_reg(366) <= "10001111101010010000011001100000";
                        f_reg(367) <= "10001100000111010000011010111000";
                        f_reg(368) <= "10001111101101110000011001100000";
                        f_reg(369) <= "00010101001101111111111111111100";
                        f_reg(370) <= "10001100000111010000011010111000";
                        f_reg(371) <= "10001111101010100000011001100100";
                        f_reg(372) <= "10001100000111010000011010111000";
                        f_reg(373) <= "10001111101110000000011001100100";
                        f_reg(374) <= "00010101010110001111111111111100";
                        f_reg(375) <= "10001100000111010000011010111000";
                        f_reg(376) <= "10001111101010110000011001101000";
                        f_reg(377) <= "10001100000111010000011010111000";
                        f_reg(378) <= "10001111101110010000011001101000";
                        f_reg(379) <= "00010101011110011111111111111100";
                        f_reg(380) <= "10001100000111010000011010111000";
                        f_reg(381) <= "10001111101011000000011001101100";
                        f_reg(382) <= "10001100000111010000011010111000";
                        f_reg(383) <= "10001111101110100000011001101100";
                        f_reg(384) <= "00010101100110101111111111111100";
                        f_reg(385) <= "10001100000111010000011010111000";
                        f_reg(386) <= "10001111101011010000011001110000";
                        f_reg(387) <= "10001100000111010000011010111000";
                        f_reg(388) <= "10001111101110110000011001110000";
                        f_reg(389) <= "00010101101110111111111111111100";
                        f_reg(390) <= "10001100000111010000011010111000";
                        f_reg(391) <= "10001111101011100000011001110100";
                        f_reg(392) <= "10001100000111010000011010111000";
                        f_reg(393) <= "10001111101111000000011001110100";
                        f_reg(394) <= "00010101110111001111111111111100";
                        f_reg(395) <= "10001100000111010000011010111000";
                        f_reg(396) <= "10001111101111100000011001111000";
                        f_reg(397) <= "10001100000111010000011010111000";
                        f_reg(398) <= "10001111101111110000011001111000";
                        f_reg(399) <= "00010111110111111111111111111100";
                        f_reg(400) <= "00010000000000001111111100110111";
                        f_reg(401) <= "00000000000000000000000000000000";
                        f_reg(402) <= "00000000000000000000000000000000";
                        f_reg(403) <= "00000000000000000000000000000000";
                        f_reg(404) <= "00000000000000000000000000000000";
                        f_reg(405) <= "00000000000000000000000000000000";
                        f_reg(406) <= "00000000000000000000000000000000";
                        f_reg(407) <= "00000000000000000000000000000000";
                        f_reg(408) <= "00000000000000000000000000000000";
                        f_reg(409) <= "00000000000000000000000000000000";
                        f_reg(410) <= "00000000000000000000000000000000";
                        f_reg(411) <= "00000000000000000000000000000000";
                        f_reg(412) <= "00000000000000000000000000000000";
                        f_reg(413) <= "00000000000000000000000000000000";
                        f_reg(414) <= "00000000000000000000000000000000";
                        f_reg(415) <= "00000000000000000000000000000000";
                        f_reg(416) <= "00000000000000000000000000000000";
                        f_reg(417) <= "00000000000000000000000000000000";
                        f_reg(418) <= "00000000000000000000000000000000";
                        f_reg(419) <= "00000000000000000000000000000000";
                        f_reg(420) <= "00000000000000000000000000000000";
                        f_reg(421) <= "00000000000000000000000000000000";
                        f_reg(422) <= "00000000000000000000000000000000";
                        f_reg(423) <= "00000000000000000000000000000000";
                        f_reg(424) <= "00000000000000000000000000000000";
                        f_reg(425) <= "00000000000000000000000000000000";
                        f_reg(426) <= "00000000000000000000000000000000";
                        f_reg(427) <= "00000000000000000000000000000000";
                        f_reg(428) <= "00000000000000000000000000000000";
                        f_reg(429) <= "00000000000000000000000000000000";
                        f_reg(430) <= "00000000000000000000000000000000";
                        f_reg(431) <= "00000000000000000000001111100111";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011000010011011111";
                        f_reg(4) <= "00101000000000100001010111011001";
                        f_reg(5) <= "00101100000000110000100011111011";
                        f_reg(6) <= "00000000010000000010000000000100";
                        f_reg(7) <= "00000000010000000010100000100011";
                        f_reg(8) <= "00000000010001010011000000100000";
                        f_reg(9) <= "00000000100001000011100000101010";
                        f_reg(10) <= "00000000111001000100000000100001";
                        f_reg(11) <= "00101100000010011011110101111111";
                        f_reg(12) <= "00000001000000000101000000100111";
                        f_reg(13) <= "00000001010010010101100000100100";
                        f_reg(14) <= "00100100111011000110110011101000";
                        f_reg(15) <= "00100000101011010111110111100101";
                        f_reg(16) <= "00101000110011100001000110000100";
                        f_reg(17) <= "00110100101011110101010110011111";
                        f_reg(18) <= "00000001000010001000000000100101";
                        f_reg(19) <= "00000001000000001000100000100010";
                        f_reg(20) <= "00000001111011011001000000100001";
                        f_reg(21) <= "00000000111000011001100000000100";
                        f_reg(22) <= "00000000101011101010000000100000";
                        f_reg(23) <= "00000010000100111010100000100000";
                        f_reg(24) <= "00000000000000000000000000000000";
                        f_reg(25) <= "00100000100101101000110010110101";
                        f_reg(26) <= "00000000000000000000000000000000";
                        f_reg(27) <= "00000010010010111011100000100010";
                        f_reg(28) <= "00000001100000001100000000100110";
                        f_reg(29) <= "00100110100110010110000001100110";
                        f_reg(30) <= "10101100000100010000001100101100";
                        f_reg(31) <= "00110010100110101011001011011010";
                        f_reg(32) <= "00000000000000000000000000000000";
                        f_reg(33) <= "10101100000110000000001100110000";
                        f_reg(34) <= "10101100000101110000001100110100";
                        f_reg(35) <= "00100110110110111010000010110001";
                        f_reg(36) <= "10101100000110100000001100111000";
                        f_reg(37) <= "00000000000000000000000000000000";
                        f_reg(38) <= "00000011011010001110000000000110";
                        f_reg(39) <= "00111100000111011101000111110000";
                        f_reg(40) <= "10101100000111000000001100111100";
                        f_reg(41) <= "00101000011111101011011110100110";
                        f_reg(42) <= "00101010110000101010010111101111";
                        f_reg(43) <= "10101100000000100000001101000000";
                        f_reg(44) <= "00111100000010100111001101000100";
                        f_reg(45) <= "00000011000111010100100000100011";
                        f_reg(46) <= "00000000000000000000000000000000";
                        f_reg(47) <= "00000011001011000011000000000110";
                        f_reg(48) <= "10101100000010000000001101000100";
                        f_reg(49) <= "00000000110101010111100000100111";
                        f_reg(50) <= "10101100000101010000001101001000";
                        f_reg(51) <= "10101100000011110000001101001100";
                        f_reg(52) <= "00000001010011010000100000101010";
                        f_reg(53) <= "00000001001111100100100000100001";
                        f_reg(54) <= "10101100000010000000001101010000";
                        f_reg(55) <= "00000000000000000000000000000000";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "00000000000000010011100011000000";
                        f_reg(58) <= "00000000000000010010101001000011";
                        f_reg(59) <= "00100001001011101100101101101010";
                        f_reg(60) <= "10101100000001110000001101010100";
                        f_reg(61) <= "10101100000001010000001101011000";
                        f_reg(62) <= "10101100000011100000001101011100";
                        f_reg(63) <= "10101100000010010000001101100000";
                        f_reg(64) <= "00100011111111111111111111111111";
                        f_reg(65) <= "00011111111000001111111111000010";
                        f_reg(66) <= "00010000000000000000000110010000";
                        f_reg(67) <= "00111100000111100000001111100111";
                        f_reg(68) <= "00111100000111110000001111100111";
                        f_reg(69) <= "00000000000111101111010000000010";
                        f_reg(70) <= "00000000000111111111110000000010";
                        f_reg(71) <= "00111100000000011000010011011111";
                        f_reg(72) <= "00111100000011111000010011011111";
                        f_reg(73) <= "00101000000000100001010111011001";
                        f_reg(74) <= "00101000000100000001010111011001";
                        f_reg(75) <= "00101100000000110000100011111011";
                        f_reg(76) <= "00101100000100010000100011111011";
                        f_reg(77) <= "00000000010000000010000000000100";
                        f_reg(78) <= "00000010000000001001000000000100";
                        f_reg(79) <= "00000000010000000010100000100011";
                        f_reg(80) <= "00000010000000001001100000100011";
                        f_reg(81) <= "00000000010001010011000000100000";
                        f_reg(82) <= "00000010000100111010000000100000";
                        f_reg(83) <= "00000000100001000011100000101010";
                        f_reg(84) <= "00000010010100101010100000101010";
                        f_reg(85) <= "00000000111001000100000000100001";
                        f_reg(86) <= "00000010101100101011000000100001";
                        f_reg(87) <= "00101100000010011011110101111111";
                        f_reg(88) <= "00101100000101111011110101111111";
                        f_reg(89) <= "00000001000000000101000000100111";
                        f_reg(90) <= "00000010110000001100000000100111";
                        f_reg(91) <= "00000001010010010101100000100100";
                        f_reg(92) <= "00000011000101111100100000100100";
                        f_reg(93) <= "00100100111011000110110011101000";
                        f_reg(94) <= "00100110101110100110110011101000";
                        f_reg(95) <= "00100000101011010111110111100101";
                        f_reg(96) <= "00100010011110110111110111100101";
                        f_reg(97) <= "00101000110011100001000110000100";
                        f_reg(98) <= "00101010100111000001000110000100";
                        f_reg(99) <= "00110100101000100101010110011111";
                        f_reg(100) <= "00110110011100000101010110011111";
                        f_reg(101) <= "00000001000010000101000000100101";
                        f_reg(102) <= "00000010110101101100000000100101";
                        f_reg(103) <= "00000001000000000100100000100010";
                        f_reg(104) <= "00000010110000001011100000100010";
                        f_reg(105) <= "00000000010011010011000000100001";
                        f_reg(106) <= "00000010000110111010000000100001";
                        f_reg(107) <= "00000000111000010001000000000100";
                        f_reg(108) <= "00000010101011111000000000000100";
                        f_reg(109) <= "00000000101011100000100000100000";
                        f_reg(110) <= "00000010011111000111100000100000";
                        f_reg(111) <= "00000001010000100011100000100000";
                        f_reg(112) <= "00000011000100001010100000100000";
                        f_reg(113) <= "00000000000000000000000000000000";
                        f_reg(114) <= "00000000000000000000000000000000";
                        f_reg(115) <= "00100000100001011000110010110101";
                        f_reg(116) <= "00100010010100111000110010110101";
                        f_reg(117) <= "00000000000000000000000000000000";
                        f_reg(118) <= "00000000000000000000000000000000";
                        f_reg(119) <= "00000000110010110111000000100010";
                        f_reg(120) <= "00000010100110011110000000100010";
                        f_reg(121) <= "00000001100000000101000000100110";
                        f_reg(122) <= "00000011010000001100000000100110";
                        f_reg(123) <= "00100100001000100110000001100110";
                        f_reg(124) <= "00100101111100000110000001100110";
                        f_reg(125) <= "00010101001101110000000011001000";
                        f_reg(126) <= "10101100000010010000001100101100";
                        f_reg(127) <= "00110000001001001011001011011010";
                        f_reg(128) <= "00110001111100101011001011011010";
                        f_reg(129) <= "00000000000000000000000000000000";
                        f_reg(130) <= "00000000000000000000000000000000";
                        f_reg(131) <= "00010101010110000000000011000010";
                        f_reg(132) <= "10101100000010100000001100110000";
                        f_reg(133) <= "00010101110111000000000011000000";
                        f_reg(134) <= "10101100000011100000001100110100";
                        f_reg(135) <= "00100100101001101010000010110001";
                        f_reg(136) <= "00100110011101001010000010110001";
                        f_reg(137) <= "00010100100100100000000010111100";
                        f_reg(138) <= "10101100000001000000001100111000";
                        f_reg(139) <= "00000000000000000000000000000000";
                        f_reg(140) <= "00000000000000000000000000000000";
                        f_reg(141) <= "00000000110010000101100000000110";
                        f_reg(142) <= "00000010100101101100100000000110";
                        f_reg(143) <= "00111100000010011101000111110000";
                        f_reg(144) <= "00111100000101111101000111110000";
                        f_reg(145) <= "00010101011110010000000010110100";
                        f_reg(146) <= "10101100000010110000001100111100";
                        f_reg(147) <= "00101000011000011011011110100110";
                        f_reg(148) <= "00101010001011111011011110100110";
                        f_reg(149) <= "00101000101011101010010111101111";
                        f_reg(150) <= "00101010011111001010010111101111";
                        f_reg(151) <= "00010101110111000000000010101110";
                        f_reg(152) <= "10101100000011100000001101000000";
                        f_reg(153) <= "00111100000001000111001101000100";
                        f_reg(154) <= "00111100000100100111001101000100";
                        f_reg(155) <= "00000001010010010011000000100011";
                        f_reg(156) <= "00000011000101111010000000100011";
                        f_reg(157) <= "00000000000000000000000000000000";
                        f_reg(158) <= "00000000000000000000000000000000";
                        f_reg(159) <= "00000000010011000101100000000110";
                        f_reg(160) <= "00000010000110101100100000000110";
                        f_reg(161) <= "00010101000101100000000010100100";
                        f_reg(162) <= "10101100000010000000001101000100";
                        f_reg(163) <= "00000001011001110001100000100111";
                        f_reg(164) <= "00000011001101011000100000100111";
                        f_reg(165) <= "00010100111101010000000010100000";
                        f_reg(166) <= "10101100000001110000001101001000";
                        f_reg(167) <= "00010100011100010000000010011110";
                        f_reg(168) <= "10101100000000110000001101001100";
                        f_reg(169) <= "00000000100011010010100000101010";
                        f_reg(170) <= "00000010010110111001100000101010";
                        f_reg(171) <= "00000000110000010011000000100001";
                        f_reg(172) <= "00000010100011111010000000100001";
                        f_reg(173) <= "00010101000101100000000010011000";
                        f_reg(174) <= "10101100000010000000001101010000";
                        f_reg(175) <= "00000000000000000000000000000000";
                        f_reg(176) <= "00000000000000000000000000000000";
                        f_reg(177) <= "00000000000000000000000000000000";
                        f_reg(178) <= "00000000000000000000000000000000";
                        f_reg(179) <= "00000000000001010111000011000000";
                        f_reg(180) <= "00000000000100111110000011000000";
                        f_reg(181) <= "00000000000001010101001001000011";
                        f_reg(182) <= "00000000000100111100001001000011";
                        f_reg(183) <= "00100000110010011100101101101010";
                        f_reg(184) <= "00100010100101111100101101101010";
                        f_reg(185) <= "00010101110111000000000010001100";
                        f_reg(186) <= "10101100000011100000001101010100";
                        f_reg(187) <= "00010101010110000000000010001010";
                        f_reg(188) <= "10101100000010100000001101011000";
                        f_reg(189) <= "00010101001101110000000010001000";
                        f_reg(190) <= "10101100000010010000001101011100";
                        f_reg(191) <= "00010100110101000000000010000110";
                        f_reg(192) <= "10101100000001100000001101100000";
                        f_reg(193) <= "00100011110111011111111100000110";
                        f_reg(194) <= "00010011101000000000000000011000";
                        f_reg(195) <= "00100011110111011111111000001100";
                        f_reg(196) <= "00010011101000000000000000010110";
                        f_reg(197) <= "00100011110111011111110100010010";
                        f_reg(198) <= "00010011101000000000000000010100";
                        f_reg(199) <= "00100011110111101111111111111111";
                        f_reg(200) <= "00100011111111111111111111111111";
                        f_reg(201) <= "00010111110111110000000001111100";
                        f_reg(202) <= "00011111111000001111111101111101";
                        f_reg(203) <= "00010000000000000000000100000111";
                        f_reg(204) <= "00000000000000000000000000000000";
                        f_reg(205) <= "00000000000000000000000000000000";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00000000000000000000000000000000";
                        f_reg(209) <= "00000000000000000000000000000000";
                        f_reg(210) <= "00000000000000000000000000000000";
                        f_reg(211) <= "00000000000000000000000000000000";
                        f_reg(212) <= "00000000000000000000000000000000";
                        f_reg(213) <= "00000000000000000000000000000000";
                        f_reg(214) <= "00000000000000000000000000000000";
                        f_reg(215) <= "00000000000000000000000000000000";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "10001100000111010000011010111000";
                        f_reg(219) <= "00011111101000000000000000000011";
                        f_reg(220) <= "00100000000111010000000000111100";
                        f_reg(221) <= "00010000000000000000000000000010";
                        f_reg(222) <= "00100000000111010000000000000000";
                        f_reg(223) <= "00010100001011110000000001100110";
                        f_reg(224) <= "10101111101000010000011001000000";
                        f_reg(225) <= "10001100000111010000011010111000";
                        f_reg(226) <= "00011111101000000000000000000011";
                        f_reg(227) <= "00100000000111010000000000111100";
                        f_reg(228) <= "00010000000000000000000000000010";
                        f_reg(229) <= "00100000000111010000000000000000";
                        f_reg(230) <= "00010100010100000000000001011111";
                        f_reg(231) <= "10101111101000100000011001000100";
                        f_reg(232) <= "10001100000111010000011010111000";
                        f_reg(233) <= "00011111101000000000000000000011";
                        f_reg(234) <= "00100000000111010000000000111100";
                        f_reg(235) <= "00010000000000000000000000000010";
                        f_reg(236) <= "00100000000111010000000000000000";
                        f_reg(237) <= "00010100011100010000000001011000";
                        f_reg(238) <= "10101111101000110000011001001000";
                        f_reg(239) <= "10001100000111010000011010111000";
                        f_reg(240) <= "00011111101000000000000000000011";
                        f_reg(241) <= "00100000000111010000000000111100";
                        f_reg(242) <= "00010000000000000000000000000010";
                        f_reg(243) <= "00100000000111010000000000000000";
                        f_reg(244) <= "00010100100100100000000001010001";
                        f_reg(245) <= "10101111101001000000011001001100";
                        f_reg(246) <= "10001100000111010000011010111000";
                        f_reg(247) <= "00011111101000000000000000000011";
                        f_reg(248) <= "00100000000111010000000000111100";
                        f_reg(249) <= "00010000000000000000000000000010";
                        f_reg(250) <= "00100000000111010000000000000000";
                        f_reg(251) <= "00010100101100110000000001001010";
                        f_reg(252) <= "10101111101001010000011001010000";
                        f_reg(253) <= "10001100000111010000011010111000";
                        f_reg(254) <= "00011111101000000000000000000011";
                        f_reg(255) <= "00100000000111010000000000111100";
                        f_reg(256) <= "00010000000000000000000000000010";
                        f_reg(257) <= "00100000000111010000000000000000";
                        f_reg(258) <= "00010100110101000000000001000011";
                        f_reg(259) <= "10101111101001100000011001010100";
                        f_reg(260) <= "10001100000111010000011010111000";
                        f_reg(261) <= "00011111101000000000000000000011";
                        f_reg(262) <= "00100000000111010000000000111100";
                        f_reg(263) <= "00010000000000000000000000000010";
                        f_reg(264) <= "00100000000111010000000000000000";
                        f_reg(265) <= "00010100111101010000000000111100";
                        f_reg(266) <= "10101111101001110000011001011000";
                        f_reg(267) <= "10001100000111010000011010111000";
                        f_reg(268) <= "00011111101000000000000000000011";
                        f_reg(269) <= "00100000000111010000000000111100";
                        f_reg(270) <= "00010000000000000000000000000010";
                        f_reg(271) <= "00100000000111010000000000000000";
                        f_reg(272) <= "00010101000101100000000000110101";
                        f_reg(273) <= "10101111101010000000011001011100";
                        f_reg(274) <= "10001100000111010000011010111000";
                        f_reg(275) <= "00011111101000000000000000000011";
                        f_reg(276) <= "00100000000111010000000000111100";
                        f_reg(277) <= "00010000000000000000000000000010";
                        f_reg(278) <= "00100000000111010000000000000000";
                        f_reg(279) <= "00010101001101110000000000101110";
                        f_reg(280) <= "10101111101010010000011001100000";
                        f_reg(281) <= "10001100000111010000011010111000";
                        f_reg(282) <= "00011111101000000000000000000011";
                        f_reg(283) <= "00100000000111010000000000111100";
                        f_reg(284) <= "00010000000000000000000000000010";
                        f_reg(285) <= "00100000000111010000000000000000";
                        f_reg(286) <= "00010101010110000000000000100111";
                        f_reg(287) <= "10101111101010100000011001100100";
                        f_reg(288) <= "10001100000111010000011010111000";
                        f_reg(289) <= "00011111101000000000000000000011";
                        f_reg(290) <= "00100000000111010000000000111100";
                        f_reg(291) <= "00010000000000000000000000000010";
                        f_reg(292) <= "00100000000111010000000000000000";
                        f_reg(293) <= "00010101011110010000000000100000";
                        f_reg(294) <= "10101111101010110000011001101000";
                        f_reg(295) <= "10001100000111010000011010111000";
                        f_reg(296) <= "00011111101000000000000000000011";
                        f_reg(297) <= "00100000000111010000000000111100";
                        f_reg(298) <= "00010000000000000000000000000010";
                        f_reg(299) <= "00100000000111010000000000000000";
                        f_reg(300) <= "00010101100110100000000000011001";
                        f_reg(301) <= "10101111101011000000011001101100";
                        f_reg(302) <= "10001100000111010000011010111000";
                        f_reg(303) <= "00011111101000000000000000000011";
                        f_reg(304) <= "00100000000111010000000000111100";
                        f_reg(305) <= "00010000000000000000000000000010";
                        f_reg(306) <= "00100000000111010000000000000000";
                        f_reg(307) <= "00010101101110110000000000010010";
                        f_reg(308) <= "10101111101011010000011001110000";
                        f_reg(309) <= "10001100000111010000011010111000";
                        f_reg(310) <= "00011111101000000000000000000011";
                        f_reg(311) <= "00100000000111010000000000111100";
                        f_reg(312) <= "00010000000000000000000000000010";
                        f_reg(313) <= "00100000000111010000000000000000";
                        f_reg(314) <= "00010101110111000000000000001011";
                        f_reg(315) <= "10101111101011100000011001110100";
                        f_reg(316) <= "10001100000111010000011010111000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010111110111110000000000000100";
                        f_reg(322) <= "10101111101111100000011001111000";
                        f_reg(323) <= "10101100000111010000011010111000";
                        f_reg(324) <= "00010000000000001111111110000011";
                        f_reg(325) <= "10001100000111010000011010111000";
                        f_reg(326) <= "10001111101000010000011001000000";
                        f_reg(327) <= "10001100000111010000011010111000";
                        f_reg(328) <= "10001111101011110000011001000000";
                        f_reg(329) <= "00010100001011111111111111111100";
                        f_reg(330) <= "10001100000111010000011010111000";
                        f_reg(331) <= "10001111101000100000011001000100";
                        f_reg(332) <= "10001100000111010000011010111000";
                        f_reg(333) <= "10001111101100000000011001000100";
                        f_reg(334) <= "00010100010100001111111111111100";
                        f_reg(335) <= "10001100000111010000011010111000";
                        f_reg(336) <= "10001111101000110000011001001000";
                        f_reg(337) <= "10001100000111010000011010111000";
                        f_reg(338) <= "10001111101100010000011001001000";
                        f_reg(339) <= "00010100011100011111111111111100";
                        f_reg(340) <= "10001100000111010000011010111000";
                        f_reg(341) <= "10001111101001000000011001001100";
                        f_reg(342) <= "10001100000111010000011010111000";
                        f_reg(343) <= "10001111101100100000011001001100";
                        f_reg(344) <= "00010100100100101111111111111100";
                        f_reg(345) <= "10001100000111010000011010111000";
                        f_reg(346) <= "10001111101001010000011001010000";
                        f_reg(347) <= "10001100000111010000011010111000";
                        f_reg(348) <= "10001111101100110000011001010000";
                        f_reg(349) <= "00010100101100111111111111111100";
                        f_reg(350) <= "10001100000111010000011010111000";
                        f_reg(351) <= "10001111101001100000011001010100";
                        f_reg(352) <= "10001100000111010000011010111000";
                        f_reg(353) <= "10001111101101000000011001010100";
                        f_reg(354) <= "00010100110101001111111111111100";
                        f_reg(355) <= "10001100000111010000011010111000";
                        f_reg(356) <= "10001111101001110000011001011000";
                        f_reg(357) <= "10001100000111010000011010111000";
                        f_reg(358) <= "10001111101101010000011001011000";
                        f_reg(359) <= "00010100111101011111111111111100";
                        f_reg(360) <= "10001100000111010000011010111000";
                        f_reg(361) <= "10001111101010000000011001011100";
                        f_reg(362) <= "10001100000111010000011010111000";
                        f_reg(363) <= "10001111101101100000011001011100";
                        f_reg(364) <= "00010101000101101111111111111100";
                        f_reg(365) <= "10001100000111010000011010111000";
                        f_reg(366) <= "10001111101010010000011001100000";
                        f_reg(367) <= "10001100000111010000011010111000";
                        f_reg(368) <= "10001111101101110000011001100000";
                        f_reg(369) <= "00010101001101111111111111111100";
                        f_reg(370) <= "10001100000111010000011010111000";
                        f_reg(371) <= "10001111101010100000011001100100";
                        f_reg(372) <= "10001100000111010000011010111000";
                        f_reg(373) <= "10001111101110000000011001100100";
                        f_reg(374) <= "00010101010110001111111111111100";
                        f_reg(375) <= "10001100000111010000011010111000";
                        f_reg(376) <= "10001111101010110000011001101000";
                        f_reg(377) <= "10001100000111010000011010111000";
                        f_reg(378) <= "10001111101110010000011001101000";
                        f_reg(379) <= "00010101011110011111111111111100";
                        f_reg(380) <= "10001100000111010000011010111000";
                        f_reg(381) <= "10001111101011000000011001101100";
                        f_reg(382) <= "10001100000111010000011010111000";
                        f_reg(383) <= "10001111101110100000011001101100";
                        f_reg(384) <= "00010101100110101111111111111100";
                        f_reg(385) <= "10001100000111010000011010111000";
                        f_reg(386) <= "10001111101011010000011001110000";
                        f_reg(387) <= "10001100000111010000011010111000";
                        f_reg(388) <= "10001111101110110000011001110000";
                        f_reg(389) <= "00010101101110111111111111111100";
                        f_reg(390) <= "10001100000111010000011010111000";
                        f_reg(391) <= "10001111101011100000011001110100";
                        f_reg(392) <= "10001100000111010000011010111000";
                        f_reg(393) <= "10001111101111000000011001110100";
                        f_reg(394) <= "00010101110111001111111111111100";
                        f_reg(395) <= "10001100000111010000011010111000";
                        f_reg(396) <= "10001111101111100000011001111000";
                        f_reg(397) <= "10001100000111010000011010111000";
                        f_reg(398) <= "10001111101111110000011001111000";
                        f_reg(399) <= "00010111110111111111111111111100";
                        f_reg(400) <= "00010000000000001111111100110111";
                        f_reg(401) <= "00000000000000000000000000000000";
                        f_reg(402) <= "00000000000000000000000000000000";
                        f_reg(403) <= "00000000000000000000000000000000";
                        f_reg(404) <= "00000000000000000000000000000000";
                        f_reg(405) <= "00000000000000000000000000000000";
                        f_reg(406) <= "00000000000000000000000000000000";
                        f_reg(407) <= "00000000000000000000000000000000";
                        f_reg(408) <= "00000000000000000000000000000000";
                        f_reg(409) <= "00000000000000000000000000000000";
                        f_reg(410) <= "00000000000000000000000000000000";
                        f_reg(411) <= "00000000000000000000000000000000";
                        f_reg(412) <= "00000000000000000000000000000000";
                        f_reg(413) <= "00000000000000000000000000000000";
                        f_reg(414) <= "00000000000000000000000000000000";
                        f_reg(415) <= "00000000000000000000000000000000";
                        f_reg(416) <= "00000000000000000000000000000000";
                        f_reg(417) <= "00000000000000000000000000000000";
                        f_reg(418) <= "00000000000000000000000000000000";
                        f_reg(419) <= "00000000000000000000000000000000";
                        f_reg(420) <= "00000000000000000000000000000000";
                        f_reg(421) <= "00000000000000000000000000000000";
                        f_reg(422) <= "00000000000000000000000000000000";
                        f_reg(423) <= "00000000000000000000000000000000";
                        f_reg(424) <= "00000000000000000000000000000000";
                        f_reg(425) <= "00000000000000000000000000000000";
                        f_reg(426) <= "00000000000000000000000000000000";
                        f_reg(427) <= "00000000000000000000000000000000";
                        f_reg(428) <= "00000000000000000000000000000000";
                        f_reg(429) <= "00000000000000000000000000000000";
                        f_reg(430) <= "00000000000000000000000000000000";
                        f_reg(431) <= "00000000000000000000001111100111";
                        f_reg(432) <= "00000000000000000000000000000000";
                        f_reg(433) <= "00000000000000000000000000000000";
                        f_reg(434) <= "00000000000000000000000000000000";
                        f_reg(435) <= "00000000000000000000000000000000";
                        f_reg(436) <= "00000000000000000000000000000000";
                        f_reg(437) <= "00000000000000000000000000000000";
                        f_reg(438) <= "00000000000000000000000000000000";
                        f_reg(439) <= "00000000000000000000000000000000";
                        f_reg(440) <= "00000000000000000000000000000000";
                        f_reg(441) <= "00000000000000000000000000000000";
                        f_reg(442) <= "00000000000000000000000000000000";
                        f_reg(443) <= "00000000000000000000000000000000";
                        f_reg(444) <= "00000000000000000000000000000000";
                        f_reg(445) <= "00000000000000000000000000000000";
                        f_reg(446) <= "00000000000000000000000000000000";
                        f_reg(447) <= "00000000000000000000000000000000";
                        f_reg(448) <= "00000000000000000000000000000000";
                        f_reg(449) <= "00000000000000000000000000000000";
                        f_reg(450) <= "00000000000000000000000000000000";
                        f_reg(451) <= "00000000000000000000000000000000";
                        f_reg(452) <= "00000000000000000000000000000000";
                        f_reg(453) <= "00000000000000000000000000000000";
                        f_reg(454) <= "00000000000000000000000000000000";
                        f_reg(455) <= "00000000000000000000000000000000";
                        f_reg(456) <= "00000000000000000000000000000000";
                        f_reg(457) <= "00000000000000000000000000000000";
                        f_reg(458) <= "00000000000000000000000000000000";
                        f_reg(459) <= "00000000000000000000000000000000";
                        f_reg(460) <= "00000000000000000000000000000000";
                        f_reg(461) <= "00000000000000000000000000000000";
                        f_reg(462) <= "00000000000000000000000000000000";
                        f_reg(463) <= "00000000000000000000000000000000";
                        f_reg(464) <= "00000000000000000000000000000000";
                        f_reg(465) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test32_Reg_COMBINED;
