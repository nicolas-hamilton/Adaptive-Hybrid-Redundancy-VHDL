--| CARRY_SELECT_ADDER_4_SC_TB
--| Tests CARRY_SELECT_ADDER_4_SC
library IEEE;
use IEEE.std_logic_1164.all;

entity CARRY_SELECT_ADDER_4_SC_TB is
end CARRY_SELECT_ADDER_4_SC_TB;

architecture testbench of CARRY_SELECT_ADDER_4_SC_TB is
	component CARRY_SELECT_ADDER_4_SC is
		port (i_A			: in  std_logic_vector(3 downto 0);
				i_B			: in  std_logic_vector(3 downto 0);
				i_C			: in  std_logic;
				o_S			: out std_logic_vector(3 downto 0);
				o_C			: out std_logic);
	end component;
	-- Declare signals
	signal w_A : std_logic_vector(3 downto 0) := (others =>'0');
	signal w_B : std_logic_vector(3 downto 0) := (others =>'0');
	signal w_C : std_logic := '0';
	signal w_S : std_logic_vector(3 downto 0);
	signal w_Cout  : std_logic;
begin
	-- Connect CARRY_SELECT_ADDER_4_SC
	u_CARRY_SELECT_ADDER_4_SC: CARRY_SELECT_ADDER_4_SC
	port map (i_A => w_A,
				 i_B => w_B,
				 i_C => w_C,
				 o_S => w_S,
				 o_C => w_Cout);
	
	-- Process for stimulating inputs		 
	stimulus: process is
	begin
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0001";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0010";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0011";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0100";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0101";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0110";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0111";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1000";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1001";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1010";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1011";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1100";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1101";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1110";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1111";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_c <= '1';
		w_B <= B"0000";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0001";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0010";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0011";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0100";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0101";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0110";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"0111";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1000";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1001";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1010";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1011";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1100";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1101";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1110";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		w_B <= B"1111";
		w_A <= B"0000";
		wait for 20 ns;
		w_A <= B"0001";
		wait for 20 ns;
		w_A <= B"0010";
		wait for 20 ns;
		w_A <= B"0011";
		wait for 20 ns;
		w_A <= B"0100";
		wait for 20 ns;
		w_A <= B"0101";
		wait for 20 ns;
		w_A <= B"0110";
		wait for 20 ns;
		w_A <= B"0111";
		wait for 20 ns;
		w_A <= B"1000";
		wait for 20 ns;
		w_A <= B"1001";
		wait for 20 ns;
		w_A <= B"1010";
		wait for 20 ns;
		w_A <= B"1011";
		wait for 20 ns;
		w_A <= B"1100";
		wait for 20 ns;
		w_A <= B"1101";
		wait for 20 ns;
		w_A <= B"1110";
		wait for 20 ns;
		w_A <= B"1111";
		wait for 20 ns;
		wait;
	end process stimulus;
end testbench;