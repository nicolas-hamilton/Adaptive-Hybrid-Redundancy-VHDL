--| Test49_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:11:23
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test49_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test49_Reg_COMBINED;

architecture a_Test49_Reg_COMBINED of Test49_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 564) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 564) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100", --  495 - 1980
      "00000000000000000000011111000000", --  496 - 1984
      "00000000000000000000011111000100", --  497 - 1988
      "00000000000000000000011111001000", --  498 - 1992
      "00000000000000000000011111001100", --  499 - 1996
      "00000000000000000000011111010000", --  500 - 2000
      "00000000000000000000011111010100", --  501 - 2004
      "00000000000000000000011111011000", --  502 - 2008
      "00000000000000000000011111011100", --  503 - 2012
      "00000000000000000000011111100000", --  504 - 2016
      "00000000000000000000011111100100", --  505 - 2020
      "00000000000000000000011111101000", --  506 - 2024
      "00000000000000000000011111101100", --  507 - 2028
      "00000000000000000000011111110000", --  508 - 2032
      "00000000000000000000011111110100", --  509 - 2036
      "00000000000000000000011111111000", --  510 - 2040
      "00000000000000000000011111111100", --  511 - 2044
      "00000000000000000000100000000000", --  512 - 2048
      "00000000000000000000100000000100", --  513 - 2052
      "00000000000000000000100000001000", --  514 - 2056
      "00000000000000000000100000001100", --  515 - 2060
      "00000000000000000000100000010000", --  516 - 2064
      "00000000000000000000100000010100", --  517 - 2068
      "00000000000000000000100000011000", --  518 - 2072
      "00000000000000000000100000011100", --  519 - 2076
      "00000000000000000000100000100000", --  520 - 2080
      "00000000000000000000100000100100", --  521 - 2084
      "00000000000000000000100000101000", --  522 - 2088
      "00000000000000000000100000101100", --  523 - 2092
      "00000000000000000000100000110000", --  524 - 2096
      "00000000000000000000100000110100", --  525 - 2100
      "00000000000000000000100000111000", --  526 - 2104
      "00000000000000000000100000111100", --  527 - 2108
      "00000000000000000000100001000000", --  528 - 2112
      "00000000000000000000100001000100", --  529 - 2116
      "00000000000000000000100001001000", --  530 - 2120
      "00000000000000000000100001001100", --  531 - 2124
      "00000000000000000000100001010000", --  532 - 2128
      "00000000000000000000100001010100", --  533 - 2132
      "00000000000000000000100001011000", --  534 - 2136
      "00000000000000000000100001011100", --  535 - 2140
      "00000000000000000000100001100000", --  536 - 2144
      "00000000000000000000100001100100", --  537 - 2148
      "00000000000000000000100001101000", --  538 - 2152
      "00000000000000000000100001101100", --  539 - 2156
      "00000000000000000000100001110000", --  540 - 2160
      "00000000000000000000100001110100", --  541 - 2164
      "00000000000000000000100001111000", --  542 - 2168
      "00000000000000000000100001111100", --  543 - 2172
      "00000000000000000000100010000000", --  544 - 2176
      "00000000000000000000100010000100", --  545 - 2180
      "00000000000000000000100010001000", --  546 - 2184
      "00000000000000000000100010001100", --  547 - 2188
      "00000000000000000000100010010000", --  548 - 2192
      "00000000000000000000100010010100", --  549 - 2196
      "00000000000000000000100010011000", --  550 - 2200
      "00000000000000000000100010011100", --  551 - 2204
      "00000000000000000000100010100000", --  552 - 2208
      "00000000000000000000100010100100", --  553 - 2212
      "00000000000000000000100010101000", --  554 - 2216
      "00000000000000000000100010101100", --  555 - 2220
      "00000000000000000000100010110000", --  556 - 2224
      "00000000000000000000100010110100", --  557 - 2228
      "00000000000000000000100010111000", --  558 - 2232
      "00000000000000000000100010111100", --  559 - 2236
      "00000000000000000000100011000000", --  560 - 2240
      "00000000000000000000100011000100", --  561 - 2244
      "00000000000000000000100011001000", --  562 - 2248
      "00000000000000000000100011001100");--  563 - 2252

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000010000111101001010", --    2 -    8
      "00111000000000101100101100111110", --    3 -   12
      "10101100000000010000010010010100", --    4 -   16
      "00000000000000000001110100000010", --    5 -   20
      "00000000001000100010000000100011", --    6 -   24
      "00111000010001010010110011000011", --    7 -   28
      "00110000100001100101101111111001", --    8 -   32
      "00000000010001100011100000100000", --    9 -   36
      "00000000011000100100000000100010", --   10 -   40
      "00100100100010011101110001100011", --   11 -   44
      "00110000011010100001111000100100", --   12 -   48
      "00000001000010000101100000000110", --   13 -   52
      "10101100000001100000010010011000", --   14 -   56
      "00000000110010010110000000100000", --   15 -   60
      "00000001001010000110100000100000", --   16 -   64
      "00000000001011000111000000000110", --   17 -   68
      "00000001110010100111100000000110", --   18 -   72
      "00101001011100000010110110100111", --   19 -   76
      "10101100000000010000010010011100", --   20 -   80
      "00000001001001001000100000000110", --   21 -   84
      "00000000001001111001000000000100", --   22 -   88
      "10101100000001100000010010100000", --   23 -   92
      "00000000000000000000000000000000", --   24 -   96
      "00000000000011001001100101000010", --   25 -  100
      "00000010010001101010000000100010", --   26 -  104
      "00000001011100001010100000100111", --   27 -  108
      "10101100000011010000010010100100", --   28 -  112
      "00000010000010011011000000100100", --   29 -  116
      "00000000100100101011100000100101", --   30 -  120
      "00000010001100111100000000100110", --   31 -  124
      "00111100000110010000101100011101", --   32 -  128
      "00000011001100111101000000100010", --   33 -  132
      "00000000000100011101100010000010", --   34 -  136
      "00000011010110101110000000000100", --   35 -  140
      "00000000000111001110100000100111", --   36 -  144
      "00101111000111101000101000001000", --   37 -  148
      "00000010110101000001000000100111", --   38 -  152
      "00000011011011110001100000100001", --   39 -  156
      "00111100000010000011100101100011", --   40 -  160
      "00000011110110010111000000100111", --   41 -  164
      "00000000000010100011101110000010", --   42 -  168
      "00000010110000000011000000100000", --   43 -  172
      "00000000000000000000000000000000", --   44 -  176
      "00100111001011011111100000101100", --   45 -  180
      "00101011110100000001110110011111", --   46 -  184
      "00000011010101010100100000100000", --   47 -  188
      "00000001011101110010000000100001", --   48 -  192
      "00000001101010011001000000100101", --   49 -  196
      "00000000111010001001100000000111", --   50 -  200
      "00000000010000111000100000100001", --   51 -  204
      "00000000000000000000000000000000", --   52 -  208
      "00101100001000010001100101111000", --   53 -  212
      "10101100000001100000010010101000", --   54 -  216
      "00000010010001011100000000100100", --   55 -  220
      "10101100000110000000010010101100", --   56 -  224
      "00000011100100001101100000100000", --   57 -  228
      "00000011011101010111100000100000", --   58 -  232
      "00000000000101010101011011000011", --   59 -  236
      "00000000100010100101000000000100", --   60 -  240
      "00000010100011001011000000101010", --   61 -  244
      "00000011101100011100100000101011", --   62 -  248
      "10101100000101010000010010110000", --   63 -  252
      "00110001010111101010010100111111", --   64 -  256
      "00000010011011101101000000000110", --   65 -  260
      "00000011001101100101100000100111", --   66 -  264
      "00100001011101111101011101010111", --   67 -  268
      "00101011110011010001110011001011", --   68 -  272
      "10101100000110100000010010110100", --   69 -  276
      "10101100000101100000010010111000", --   70 -  280
      "10101100000011110000010010111100", --   71 -  284
      "10101100000110100000010011000000", --   72 -  288
      "00111011001010011011111110101011", --   73 -  292
      "00101010111010001011000111001110", --   74 -  296
      "10101100000000010000010011000100", --   75 -  300
      "10101100000010000000010011001000", --   76 -  304
      "00100001001001110011010101111100", --   77 -  308
      "10101100000100110000010011001100", --   78 -  312
      "00000000111101110001000000100100", --   79 -  316
      "00100000010000110001001001100010", --   80 -  320
      "10101100000011010000010011010000", --   81 -  324
      "10101100000000110000010011010100", --   82 -  328
      "00100011111111111111111111111111", --   83 -  332
      "00011111111000001111111110101110", --   84 -  336
      "00010000000000000000000111011110", --   85 -  340
      "00111100000111100000001111100111", --   86 -  344
      "00111100000111110000001111100111", --   87 -  348
      "00000000000111101111010000000010", --   88 -  352
      "00000000000111111111110000000010", --   89 -  356
      "00111100000000010000111101001010", --   90 -  360
      "00111100000011110000111101001010", --   91 -  364
      "00111000000000101100101100111110", --   92 -  368
      "00111000000100001100101100111110", --   93 -  372
      "00010100001011110000000101001000", --   94 -  376
      "10101100000000010000010010010100", --   95 -  380
      "00000000000000000001110100000010", --   96 -  384
      "00000000000000001000110100000010", --   97 -  388
      "00000000001000100010000000100011", --   98 -  392
      "00000001111100001001000000100011", --   99 -  396
      "00111000010001010010110011000011", --  100 -  400
      "00111010000100110010110011000011", --  101 -  404
      "00110000100001100101101111111001", --  102 -  408
      "00110010010101000101101111111001", --  103 -  412
      "00000000010001100011100000100000", --  104 -  416
      "00000010000101001010100000100000", --  105 -  420
      "00000000011000100100000000100010", --  106 -  424
      "00000010001100001011000000100010", --  107 -  428
      "00100100100010011101110001100011", --  108 -  432
      "00100110010101111101110001100011", --  109 -  436
      "00110000011010100001111000100100", --  110 -  440
      "00110010001110000001111000100100", --  111 -  444
      "00000001000010000101100000000110", --  112 -  448
      "00000010110101101100100000000110", --  113 -  452
      "00010100110101000000000100110100", --  114 -  456
      "10101100000001100000010010011000", --  115 -  460
      "00000000110010010110000000100000", --  116 -  464
      "00000010100101111101000000100000", --  117 -  468
      "00000001001010000110100000100000", --  118 -  472
      "00000010111101101101100000100000", --  119 -  476
      "00000000001011000111000000000110", --  120 -  480
      "00000001111110101110000000000110", --  121 -  484
      "00000001110010100001000000000110", --  122 -  488
      "00000011100110001000000000000110", --  123 -  492
      "00101001011000110010110110100111", --  124 -  496
      "00101011001100010010110110100111", --  125 -  500
      "00010100001011110000000100101000", --  126 -  504
      "10101100000000010000010010011100", --  127 -  508
      "00000001001001000100000000000110", --  128 -  512
      "00000010111100101011000000000110", --  129 -  516
      "00000000001001110111000000000100", --  130 -  520
      "00000001111101011110000000000100", --  131 -  524
      "00010100110101000000000100100010", --  132 -  528
      "10101100000001100000010010100000", --  133 -  532
      "00000000000000000000000000000000", --  134 -  536
      "00000000000000000000000000000000", --  135 -  540
      "00000000000011000011100101000010", --  136 -  544
      "00000000000110101010100101000010", --  137 -  548
      "00010101100110100000000100011100", --  138 -  552
      "10101100000011000000010011011000", --  139 -  556
      "00000001110001100110000000100010", --  140 -  560
      "00000011100101001101000000100010", --  141 -  564
      "00000001011000110011000000100111", --  142 -  568
      "00000011001100011010000000100111", --  143 -  572
      "00010101101110110000000100010110", --  144 -  576
      "10101100000011010000010010100100", --  145 -  580
      "00000000011010010110100000100100", --  146 -  584
      "00000010001101111101100000100100", --  147 -  588
      "00000000100011100001100000100101", --  148 -  592
      "00000010010111001000100000100101", --  149 -  596
      "00000001000001110100100000100110", --  150 -  600
      "00000010110101011011100000100110", --  151 -  604
      "00111100000001000000101100011101", --  152 -  608
      "00111100000100100000101100011101", --  153 -  612
      "00000000100001110111000000100010", --  154 -  616
      "00000010010101011110000000100010", --  155 -  620
      "00000000000010000011100010000010", --  156 -  624
      "00000000000101101010100010000010", --  157 -  628
      "00000001110011100100000000000100", --  158 -  632
      "00000011100111001011000000000100", --  159 -  636
      "00010100110101000000000100000110", --  160 -  640
      "10101100000001100000010011011100", --  161 -  644
      "00000000000010000011000000100111", --  162 -  648
      "00000000000101101010000000100111", --  163 -  652
      "00010100110101000000000100000010", --  164 -  656
      "10101100000001100000010011100000", --  165 -  660
      "00101101001001101000101000001000", --  166 -  664
      "00101110111101001000101000001000", --  167 -  668
      "00000001101011000100100000100111", --  168 -  672
      "00000011011110101011100000100111", --  169 -  676
      "00010101100110100000000011111100", --  170 -  680
      "10101100000011000000010011100100", --  171 -  684
      "00000000111000100110000000100001", --  172 -  688
      "00000010101100001101000000100001", --  173 -  692
      "00111100000001110011100101100011", --  174 -  696
      "00111100000101010011100101100011", --  175 -  700
      "00000000110001000001000000100111", --  176 -  704
      "00000010100100101000000000100111", --  177 -  708
      "00010100010100000000000011110100", --  178 -  712
      "10101100000000100000010011101000", --  179 -  716
      "00000000000010100001001110000010", --  180 -  720
      "00000000000110001000001110000010", --  181 -  724
      "00000001101000000101000000100000", --  182 -  728
      "00000011011000001100000000100000", --  183 -  732
      "00000000000000000000000000000000", --  184 -  736
      "00000000000000000000000000000000", --  185 -  740
      "00100100100011011111100000101100", --  186 -  744
      "00100110010110111111100000101100", --  187 -  748
      "00101000110001000001110110011111", --  188 -  752
      "00101010100100100001110110011111", --  189 -  756
      "10001100000001100000010011011100", --  190 -  760
      "10001100000101000000010011011100", --  191 -  764
      "00010100110101001111111111111110", --  192 -  768
      "00010101000101100000000011100101", --  193 -  772
      "10101100000010000000010011011100", --  194 -  776
      "00000001110001100100000000100000", --  195 -  780
      "00000011100101001011000000100000", --  196 -  784
      "00000001011000110111000000100001", --  197 -  788
      "00000011001100011110000000100001", --  198 -  792
      "00000001101010000101100000100101", --  199 -  796
      "00000011011101101100100000100101", --  200 -  800
      "00000000010001110001100000000111", --  201 -  804
      "00000010000101011000100000000111", --  202 -  808
      "00000001001011000110100000100001", --  203 -  812
      "00000010111110101101100000100001", --  204 -  816
      "00000000000000000000000000000000", --  205 -  820
      "00000000000000000000000000000000", --  206 -  824
      "00101100001000010001100101111000", --  207 -  828
      "00101101111011110001100101111000", --  208 -  832
      "00010101010110000000000011010101", --  209 -  836
      "10101100000010100000010010101000", --  210 -  840
      "00000001011001010100000000100100", --  211 -  844
      "00000011001100111011000000100100", --  212 -  848
      "00010101000101100000000011010001", --  213 -  852
      "10101100000010000000010010101100", --  214 -  856
      "10001100000001110000010011011100", --  215 -  860
      "10001100000101010000010011011100", --  216 -  864
      "00010100111101011111111111111110", --  217 -  868
      "00000000111001000001000000100000", --  218 -  872
      "00000010101100101000000000100000", --  219 -  876
      "00000000010001100100100000100000", --  220 -  880
      "00000010000101001011100000100000", --  221 -  884
      "00000000000001100110011011000011", --  222 -  888
      "00000000000101001101011011000011", --  223 -  892
      "00000001110011000110000000000100", --  224 -  896
      "00000011100110101101000000000100", --  225 -  900
      "10001100000010100000010011100100", --  226 -  904
      "10001100000110000000010011100100", --  227 -  908
      "00010101010110001111111111111110", --  228 -  912
      "10001100000010110000010011011000", --  229 -  916
      "10001100000110010000010011011000", --  230 -  920
      "00010101011110011111111111111110", --  231 -  924
      "00000001010010110010100000101010", --  232 -  928
      "00000011000110011001100000101010", --  233 -  932
      "10001100000010000000010011100000", --  234 -  936
      "10001100000101100000010011100000", --  235 -  940
      "00010101000101101111111111111110", --  236 -  944
      "00000001000011010011100000101011", --  237 -  948
      "00000010110110111010100000101011", --  238 -  952
      "00010100110101000000000010110111", --  239 -  956
      "10101100000001100000010010110000", --  240 -  960
      "00110001100001001010010100111111", --  241 -  964
      "00110011010100101010010100111111", --  242 -  968
      "10001100000000100000010011101000", --  243 -  972
      "10001100000100000000010011101000", --  244 -  976
      "00010100010100001111111111111110", --  245 -  980
      "00000000011000100111000000000110", --  246 -  984
      "00000010001100001110000000000110", --  247 -  988
      "00000000111001010101000000100111", --  248 -  992
      "00000010101100111100000000100111", --  249 -  996
      "00100001010010111101011101010111", --  250 - 1000
      "00100011000110011101011101010111", --  251 - 1004
      "00101000100010000001110011001011", --  252 - 1008
      "00101010010101100001110011001011", --  253 - 1012
      "00010101110111000000000010101000", --  254 - 1016
      "10101100000011100000010010110100", --  255 - 1020
      "00010100101100110000000010100110", --  256 - 1024
      "10101100000001010000010010111000", --  257 - 1028
      "00010101001101110000000010100100", --  258 - 1032
      "10101100000010010000010010111100", --  259 - 1036
      "00010101110111000000000010100010", --  260 - 1040
      "10101100000011100000010011000000", --  261 - 1044
      "00111000111011011011111110101011", --  262 - 1048
      "00111010101110111011111110101011", --  263 - 1052
      "00101001011001101011000111001110", --  264 - 1056
      "00101011001101001011000111001110", --  265 - 1060
      "00010100001011110000000010011100", --  266 - 1064
      "10101100000000010000010011000100", --  267 - 1068
      "00010100110101000000000010011010", --  268 - 1072
      "10101100000001100000010011001000", --  269 - 1076
      "00100001101011000011010101111100", --  270 - 1080
      "00100011011110100011010101111100", --  271 - 1084
      "00010100011100010000000010010110", --  272 - 1088
      "10101100000000110000010011001100", --  273 - 1092
      "00000001100010110001000000100100", --  274 - 1096
      "00000011010110011000000000100100", --  275 - 1100
      "00100000010010100001001001100010", --  276 - 1104
      "00100010000110000001001001100010", --  277 - 1108
      "00010101000101100000000010010000", --  278 - 1112
      "10101100000010000000010011010000", --  279 - 1116
      "00010101010110000000000010001110", --  280 - 1120
      "10101100000010100000010011010100", --  281 - 1124
      "00100011110111011111111100000110", --  282 - 1128
      "00010011101000000000000000100000", --  283 - 1132
      "00100011110111011111111000001100", --  284 - 1136
      "00010011101000000000000000011110", --  285 - 1140
      "00100011110111011111110100010010", --  286 - 1144
      "00010011101000000000000000011100", --  287 - 1148
      "00100011110111101111111111111111", --  288 - 1152
      "00100011111111111111111111111111", --  289 - 1156
      "00010111110111110000000010000100", --  290 - 1160
      "00011111111000001111111100110111", --  291 - 1164
      "00010000000000000000000100001111", --  292 - 1168
      "00000000000000000000000000000000", --  293 - 1172
      "00000000000000000000000000000000", --  294 - 1176
      "00000000000000000000000000000000", --  295 - 1180
      "00000000000000000000000000000000", --  296 - 1184
      "00000000000000000000000000000000", --  297 - 1188
      "00000000000000000000000000000000", --  298 - 1192
      "00000000000000000000000000000000", --  299 - 1196
      "00000000000000000000000000000000", --  300 - 1200
      "00000000000000000000000000000000", --  301 - 1204
      "00000000000000000000000000000000", --  302 - 1208
      "00000000000000000000000000000000", --  303 - 1212
      "00000000000000000000000000000000", --  304 - 1216
      "00000000000000000000000000000000", --  305 - 1220
      "00000000000000000000000000000000", --  306 - 1224
      "00000000000000000000000000000000", --  307 - 1228
      "00000000000000000000000000000000", --  308 - 1232
      "00000000000000000000000000000000", --  309 - 1236
      "00000000000000000000000000000000", --  310 - 1240
      "00000000000000000000000000000000", --  311 - 1244
      "00000000000000000000000000000000", --  312 - 1248
      "00000000000000000000000000000000", --  313 - 1252
      "00000000000000000000000000000000", --  314 - 1256
      "10001100000111010000100001000000", --  315 - 1260
      "00011111101000000000000000000011", --  316 - 1264
      "00100000000111010000000000111100", --  317 - 1268
      "00010000000000000000000000000010", --  318 - 1272
      "00100000000111010000000000000000", --  319 - 1276
      "00010100001011110000000001100110", --  320 - 1280
      "10101111101000010000011111001000", --  321 - 1284
      "10001100000111010000100001000000", --  322 - 1288
      "00011111101000000000000000000011", --  323 - 1292
      "00100000000111010000000000111100", --  324 - 1296
      "00010000000000000000000000000010", --  325 - 1300
      "00100000000111010000000000000000", --  326 - 1304
      "00010100010100000000000001011111", --  327 - 1308
      "10101111101000100000011111001100", --  328 - 1312
      "10001100000111010000100001000000", --  329 - 1316
      "00011111101000000000000000000011", --  330 - 1320
      "00100000000111010000000000111100", --  331 - 1324
      "00010000000000000000000000000010", --  332 - 1328
      "00100000000111010000000000000000", --  333 - 1332
      "00010100011100010000000001011000", --  334 - 1336
      "10101111101000110000011111010000", --  335 - 1340
      "10001100000111010000100001000000", --  336 - 1344
      "00011111101000000000000000000011", --  337 - 1348
      "00100000000111010000000000111100", --  338 - 1352
      "00010000000000000000000000000010", --  339 - 1356
      "00100000000111010000000000000000", --  340 - 1360
      "00010100100100100000000001010001", --  341 - 1364
      "10101111101001000000011111010100", --  342 - 1368
      "10001100000111010000100001000000", --  343 - 1372
      "00011111101000000000000000000011", --  344 - 1376
      "00100000000111010000000000111100", --  345 - 1380
      "00010000000000000000000000000010", --  346 - 1384
      "00100000000111010000000000000000", --  347 - 1388
      "00010100101100110000000001001010", --  348 - 1392
      "10101111101001010000011111011000", --  349 - 1396
      "10001100000111010000100001000000", --  350 - 1400
      "00011111101000000000000000000011", --  351 - 1404
      "00100000000111010000000000111100", --  352 - 1408
      "00010000000000000000000000000010", --  353 - 1412
      "00100000000111010000000000000000", --  354 - 1416
      "00010100110101000000000001000011", --  355 - 1420
      "10101111101001100000011111011100", --  356 - 1424
      "10001100000111010000100001000000", --  357 - 1428
      "00011111101000000000000000000011", --  358 - 1432
      "00100000000111010000000000111100", --  359 - 1436
      "00010000000000000000000000000010", --  360 - 1440
      "00100000000111010000000000000000", --  361 - 1444
      "00010100111101010000000000111100", --  362 - 1448
      "10101111101001110000011111100000", --  363 - 1452
      "10001100000111010000100001000000", --  364 - 1456
      "00011111101000000000000000000011", --  365 - 1460
      "00100000000111010000000000111100", --  366 - 1464
      "00010000000000000000000000000010", --  367 - 1468
      "00100000000111010000000000000000", --  368 - 1472
      "00010101000101100000000000110101", --  369 - 1476
      "10101111101010000000011111100100", --  370 - 1480
      "10001100000111010000100001000000", --  371 - 1484
      "00011111101000000000000000000011", --  372 - 1488
      "00100000000111010000000000111100", --  373 - 1492
      "00010000000000000000000000000010", --  374 - 1496
      "00100000000111010000000000000000", --  375 - 1500
      "00010101001101110000000000101110", --  376 - 1504
      "10101111101010010000011111101000", --  377 - 1508
      "10001100000111010000100001000000", --  378 - 1512
      "00011111101000000000000000000011", --  379 - 1516
      "00100000000111010000000000111100", --  380 - 1520
      "00010000000000000000000000000010", --  381 - 1524
      "00100000000111010000000000000000", --  382 - 1528
      "00010101010110000000000000100111", --  383 - 1532
      "10101111101010100000011111101100", --  384 - 1536
      "10001100000111010000100001000000", --  385 - 1540
      "00011111101000000000000000000011", --  386 - 1544
      "00100000000111010000000000111100", --  387 - 1548
      "00010000000000000000000000000010", --  388 - 1552
      "00100000000111010000000000000000", --  389 - 1556
      "00010101011110010000000000100000", --  390 - 1560
      "10101111101010110000011111110000", --  391 - 1564
      "10001100000111010000100001000000", --  392 - 1568
      "00011111101000000000000000000011", --  393 - 1572
      "00100000000111010000000000111100", --  394 - 1576
      "00010000000000000000000000000010", --  395 - 1580
      "00100000000111010000000000000000", --  396 - 1584
      "00010101100110100000000000011001", --  397 - 1588
      "10101111101011000000011111110100", --  398 - 1592
      "10001100000111010000100001000000", --  399 - 1596
      "00011111101000000000000000000011", --  400 - 1600
      "00100000000111010000000000111100", --  401 - 1604
      "00010000000000000000000000000010", --  402 - 1608
      "00100000000111010000000000000000", --  403 - 1612
      "00010101101110110000000000010010", --  404 - 1616
      "10101111101011010000011111111000", --  405 - 1620
      "10001100000111010000100001000000", --  406 - 1624
      "00011111101000000000000000000011", --  407 - 1628
      "00100000000111010000000000111100", --  408 - 1632
      "00010000000000000000000000000010", --  409 - 1636
      "00100000000111010000000000000000", --  410 - 1640
      "00010101110111000000000000001011", --  411 - 1644
      "10101111101011100000011111111100", --  412 - 1648
      "10001100000111010000100001000000", --  413 - 1652
      "00011111101000000000000000000011", --  414 - 1656
      "00100000000111010000000000111100", --  415 - 1660
      "00010000000000000000000000000010", --  416 - 1664
      "00100000000111010000000000000000", --  417 - 1668
      "00010111110111110000000000000100", --  418 - 1672
      "10101111101111100000100000000000", --  419 - 1676
      "10101100000111010000100001000000", --  420 - 1680
      "00010000000000001111111101111011", --  421 - 1684
      "10001100000111010000100001000000", --  422 - 1688
      "10001111101000010000011111001000", --  423 - 1692
      "10001100000111010000100001000000", --  424 - 1696
      "10001111101011110000011111001000", --  425 - 1700
      "00010100001011111111111111111100", --  426 - 1704
      "10001100000111010000100001000000", --  427 - 1708
      "10001111101000100000011111001100", --  428 - 1712
      "10001100000111010000100001000000", --  429 - 1716
      "10001111101100000000011111001100", --  430 - 1720
      "00010100010100001111111111111100", --  431 - 1724
      "10001100000111010000100001000000", --  432 - 1728
      "10001111101000110000011111010000", --  433 - 1732
      "10001100000111010000100001000000", --  434 - 1736
      "10001111101100010000011111010000", --  435 - 1740
      "00010100011100011111111111111100", --  436 - 1744
      "10001100000111010000100001000000", --  437 - 1748
      "10001111101001000000011111010100", --  438 - 1752
      "10001100000111010000100001000000", --  439 - 1756
      "10001111101100100000011111010100", --  440 - 1760
      "00010100100100101111111111111100", --  441 - 1764
      "10001100000111010000100001000000", --  442 - 1768
      "10001111101001010000011111011000", --  443 - 1772
      "10001100000111010000100001000000", --  444 - 1776
      "10001111101100110000011111011000", --  445 - 1780
      "00010100101100111111111111111100", --  446 - 1784
      "10001100000111010000100001000000", --  447 - 1788
      "10001111101001100000011111011100", --  448 - 1792
      "10001100000111010000100001000000", --  449 - 1796
      "10001111101101000000011111011100", --  450 - 1800
      "00010100110101001111111111111100", --  451 - 1804
      "10001100000111010000100001000000", --  452 - 1808
      "10001111101001110000011111100000", --  453 - 1812
      "10001100000111010000100001000000", --  454 - 1816
      "10001111101101010000011111100000", --  455 - 1820
      "00010100111101011111111111111100", --  456 - 1824
      "10001100000111010000100001000000", --  457 - 1828
      "10001111101010000000011111100100", --  458 - 1832
      "10001100000111010000100001000000", --  459 - 1836
      "10001111101101100000011111100100", --  460 - 1840
      "00010101000101101111111111111100", --  461 - 1844
      "10001100000111010000100001000000", --  462 - 1848
      "10001111101010010000011111101000", --  463 - 1852
      "10001100000111010000100001000000", --  464 - 1856
      "10001111101101110000011111101000", --  465 - 1860
      "00010101001101111111111111111100", --  466 - 1864
      "10001100000111010000100001000000", --  467 - 1868
      "10001111101010100000011111101100", --  468 - 1872
      "10001100000111010000100001000000", --  469 - 1876
      "10001111101110000000011111101100", --  470 - 1880
      "00010101010110001111111111111100", --  471 - 1884
      "10001100000111010000100001000000", --  472 - 1888
      "10001111101010110000011111110000", --  473 - 1892
      "10001100000111010000100001000000", --  474 - 1896
      "10001111101110010000011111110000", --  475 - 1900
      "00010101011110011111111111111100", --  476 - 1904
      "10001100000111010000100001000000", --  477 - 1908
      "10001111101011000000011111110100", --  478 - 1912
      "10001100000111010000100001000000", --  479 - 1916
      "10001111101110100000011111110100", --  480 - 1920
      "00010101100110101111111111111100", --  481 - 1924
      "10001100000111010000100001000000", --  482 - 1928
      "10001111101011010000011111111000", --  483 - 1932
      "10001100000111010000100001000000", --  484 - 1936
      "10001111101110110000011111111000", --  485 - 1940
      "00010101101110111111111111111100", --  486 - 1944
      "10001100000111010000100001000000", --  487 - 1948
      "10001111101011100000011111111100", --  488 - 1952
      "10001100000111010000100001000000", --  489 - 1956
      "10001111101111000000011111111100", --  490 - 1960
      "00010101110111001111111111111100", --  491 - 1964
      "10001100000111010000100001000000", --  492 - 1968
      "10001111101111100000100000000000", --  493 - 1972
      "10001100000111010000100001000000", --  494 - 1976
      "10001111101111110000100000000000", --  495 - 1980
      "00010111110111111111111111111100", --  496 - 1984
      "00010000000000001111111100101111", --  497 - 1988
      "00000000000000000000000000000000", --  498 - 1992
      "00000000000000000000000000000000", --  499 - 1996
      "00000000000000000000000000000000", --  500 - 2000
      "00000000000000000000000000000000", --  501 - 2004
      "00000000000000000000000000000000", --  502 - 2008
      "00000000000000000000000000000000", --  503 - 2012
      "00000000000000000000000000000000", --  504 - 2016
      "00000000000000000000000000000000", --  505 - 2020
      "00000000000000000000000000000000", --  506 - 2024
      "00000000000000000000000000000000", --  507 - 2028
      "00000000000000000000000000000000", --  508 - 2032
      "00000000000000000000000000000000", --  509 - 2036
      "00000000000000000000000000000000", --  510 - 2040
      "00000000000000000000000000000000", --  511 - 2044
      "00000000000000000000000000000000", --  512 - 2048
      "00000000000000000000000000000000", --  513 - 2052
      "00000000000000000000000000000000", --  514 - 2056
      "00000000000000000000000000000000", --  515 - 2060
      "00000000000000000000000000000000", --  516 - 2064
      "00000000000000000000000000000000", --  517 - 2068
      "00000000000000000000000000000000", --  518 - 2072
      "00000000000000000000000000000000", --  519 - 2076
      "00000000000000000000000000000000", --  520 - 2080
      "00000000000000000000000000000000", --  521 - 2084
      "00000000000000000000000000000000", --  522 - 2088
      "00000000000000000000000000000000", --  523 - 2092
      "00000000000000000000000000000000", --  524 - 2096
      "00000000000000000000000000000000", --  525 - 2100
      "00000000000000000000000000000000", --  526 - 2104
      "00000000000000000000000000000000", --  527 - 2108
      "00000000000000000000001111100111", --  528 - 2112
      "00000000000000000000000000000000", --  529 - 2116
      "00000000000000000000000000000000", --  530 - 2120
      "00000000000000000000000000000000", --  531 - 2124
      "00000000000000000000000000000000", --  532 - 2128
      "00000000000000000000000000000000", --  533 - 2132
      "00000000000000000000000000000000", --  534 - 2136
      "00000000000000000000000000000000", --  535 - 2140
      "00000000000000000000000000000000", --  536 - 2144
      "00000000000000000000000000000000", --  537 - 2148
      "00000000000000000000000000000000", --  538 - 2152
      "00000000000000000000000000000000", --  539 - 2156
      "00000000000000000000000000000000", --  540 - 2160
      "00000000000000000000000000000000", --  541 - 2164
      "00000000000000000000000000000000", --  542 - 2168
      "00000000000000000000000000000000", --  543 - 2172
      "00000000000000000000000000000000", --  544 - 2176
      "00000000000000000000000000000000", --  545 - 2180
      "00000000000000000000000000000000", --  546 - 2184
      "00000000000000000000000000000000", --  547 - 2188
      "00000000000000000000000000000000", --  548 - 2192
      "00000000000000000000000000000000", --  549 - 2196
      "00000000000000000000000000000000", --  550 - 2200
      "00000000000000000000000000000000", --  551 - 2204
      "00000000000000000000000000000000", --  552 - 2208
      "00000000000000000000000000000000", --  553 - 2212
      "00000000000000000000000000000000", --  554 - 2216
      "00000000000000000000000000000000", --  555 - 2220
      "00000000000000000000000000000000", --  556 - 2224
      "00000000000000000000000000000000", --  557 - 2228
      "00000000000000000000000000000000", --  558 - 2232
      "00000000000000000000000000000000", --  559 - 2236
      "00000000000000000000000000000000", --  560 - 2240
      "00000000000000000000000000000000", --  561 - 2244
      "00000000000000000000000000000000", --  562 - 2248
      "00000000000000000000000000000000");--  563 - 2252

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000010000111101001010";
         f_reg(4) <= "00111000000000101100101100111110";
         f_reg(5) <= "10101100000000010000010010010100";
         f_reg(6) <= "00000000000000000001110100000010";
         f_reg(7) <= "00000000001000100010000000100011";
         f_reg(8) <= "00111000010001010010110011000011";
         f_reg(9) <= "00110000100001100101101111111001";
         f_reg(10) <= "00000000010001100011100000100000";
         f_reg(11) <= "00000000011000100100000000100010";
         f_reg(12) <= "00100100100010011101110001100011";
         f_reg(13) <= "00110000011010100001111000100100";
         f_reg(14) <= "00000001000010000101100000000110";
         f_reg(15) <= "10101100000001100000010010011000";
         f_reg(16) <= "00000000110010010110000000100000";
         f_reg(17) <= "00000001001010000110100000100000";
         f_reg(18) <= "00000000001011000111000000000110";
         f_reg(19) <= "00000001110010100111100000000110";
         f_reg(20) <= "00101001011100000010110110100111";
         f_reg(21) <= "10101100000000010000010010011100";
         f_reg(22) <= "00000001001001001000100000000110";
         f_reg(23) <= "00000000001001111001000000000100";
         f_reg(24) <= "10101100000001100000010010100000";
         f_reg(25) <= "00000000000000000000000000000000";
         f_reg(26) <= "00000000000011001001100101000010";
         f_reg(27) <= "00000010010001101010000000100010";
         f_reg(28) <= "00000001011100001010100000100111";
         f_reg(29) <= "10101100000011010000010010100100";
         f_reg(30) <= "00000010000010011011000000100100";
         f_reg(31) <= "00000000100100101011100000100101";
         f_reg(32) <= "00000010001100111100000000100110";
         f_reg(33) <= "00111100000110010000101100011101";
         f_reg(34) <= "00000011001100111101000000100010";
         f_reg(35) <= "00000000000100011101100010000010";
         f_reg(36) <= "00000011010110101110000000000100";
         f_reg(37) <= "00000000000111001110100000100111";
         f_reg(38) <= "00101111000111101000101000001000";
         f_reg(39) <= "00000010110101000001000000100111";
         f_reg(40) <= "00000011011011110001100000100001";
         f_reg(41) <= "00111100000010000011100101100011";
         f_reg(42) <= "00000011110110010111000000100111";
         f_reg(43) <= "00000000000010100011101110000010";
         f_reg(44) <= "00000010110000000011000000100000";
         f_reg(45) <= "00000000000000000000000000000000";
         f_reg(46) <= "00100111001011011111100000101100";
         f_reg(47) <= "00101011110100000001110110011111";
         f_reg(48) <= "00000011010101010100100000100000";
         f_reg(49) <= "00000001011101110010000000100001";
         f_reg(50) <= "00000001101010011001000000100101";
         f_reg(51) <= "00000000111010001001100000000111";
         f_reg(52) <= "00000000010000111000100000100001";
         f_reg(53) <= "00000000000000000000000000000000";
         f_reg(54) <= "00101100001000010001100101111000";
         f_reg(55) <= "10101100000001100000010010101000";
         f_reg(56) <= "00000010010001011100000000100100";
         f_reg(57) <= "10101100000110000000010010101100";
         f_reg(58) <= "00000011100100001101100000100000";
         f_reg(59) <= "00000011011101010111100000100000";
         f_reg(60) <= "00000000000101010101011011000011";
         f_reg(61) <= "00000000100010100101000000000100";
         f_reg(62) <= "00000010100011001011000000101010";
         f_reg(63) <= "00000011101100011100100000101011";
         f_reg(64) <= "10101100000101010000010010110000";
         f_reg(65) <= "00110001010111101010010100111111";
         f_reg(66) <= "00000010011011101101000000000110";
         f_reg(67) <= "00000011001101100101100000100111";
         f_reg(68) <= "00100001011101111101011101010111";
         f_reg(69) <= "00101011110011010001110011001011";
         f_reg(70) <= "10101100000110100000010010110100";
         f_reg(71) <= "10101100000101100000010010111000";
         f_reg(72) <= "10101100000011110000010010111100";
         f_reg(73) <= "10101100000110100000010011000000";
         f_reg(74) <= "00111011001010011011111110101011";
         f_reg(75) <= "00101010111010001011000111001110";
         f_reg(76) <= "10101100000000010000010011000100";
         f_reg(77) <= "10101100000010000000010011001000";
         f_reg(78) <= "00100001001001110011010101111100";
         f_reg(79) <= "10101100000100110000010011001100";
         f_reg(80) <= "00000000111101110001000000100100";
         f_reg(81) <= "00100000010000110001001001100010";
         f_reg(82) <= "10101100000011010000010011010000";
         f_reg(83) <= "10101100000000110000010011010100";
         f_reg(84) <= "00100011111111111111111111111111";
         f_reg(85) <= "00011111111000001111111110101110";
         f_reg(86) <= "00010000000000000000000111011110";
         f_reg(87) <= "00111100000111100000001111100111";
         f_reg(88) <= "00111100000111110000001111100111";
         f_reg(89) <= "00000000000111101111010000000010";
         f_reg(90) <= "00000000000111111111110000000010";
         f_reg(91) <= "00111100000000010000111101001010";
         f_reg(92) <= "00111100000011110000111101001010";
         f_reg(93) <= "00111000000000101100101100111110";
         f_reg(94) <= "00111000000100001100101100111110";
         f_reg(95) <= "00010100001011110000000101001000";
         f_reg(96) <= "10101100000000010000010010010100";
         f_reg(97) <= "00000000000000000001110100000010";
         f_reg(98) <= "00000000000000001000110100000010";
         f_reg(99) <= "00000000001000100010000000100011";
         f_reg(100) <= "00000001111100001001000000100011";
         f_reg(101) <= "00111000010001010010110011000011";
         f_reg(102) <= "00111010000100110010110011000011";
         f_reg(103) <= "00110000100001100101101111111001";
         f_reg(104) <= "00110010010101000101101111111001";
         f_reg(105) <= "00000000010001100011100000100000";
         f_reg(106) <= "00000010000101001010100000100000";
         f_reg(107) <= "00000000011000100100000000100010";
         f_reg(108) <= "00000010001100001011000000100010";
         f_reg(109) <= "00100100100010011101110001100011";
         f_reg(110) <= "00100110010101111101110001100011";
         f_reg(111) <= "00110000011010100001111000100100";
         f_reg(112) <= "00110010001110000001111000100100";
         f_reg(113) <= "00000001000010000101100000000110";
         f_reg(114) <= "00000010110101101100100000000110";
         f_reg(115) <= "00010100110101000000000100110100";
         f_reg(116) <= "10101100000001100000010010011000";
         f_reg(117) <= "00000000110010010110000000100000";
         f_reg(118) <= "00000010100101111101000000100000";
         f_reg(119) <= "00000001001010000110100000100000";
         f_reg(120) <= "00000010111101101101100000100000";
         f_reg(121) <= "00000000001011000111000000000110";
         f_reg(122) <= "00000001111110101110000000000110";
         f_reg(123) <= "00000001110010100001000000000110";
         f_reg(124) <= "00000011100110001000000000000110";
         f_reg(125) <= "00101001011000110010110110100111";
         f_reg(126) <= "00101011001100010010110110100111";
         f_reg(127) <= "00010100001011110000000100101000";
         f_reg(128) <= "10101100000000010000010010011100";
         f_reg(129) <= "00000001001001000100000000000110";
         f_reg(130) <= "00000010111100101011000000000110";
         f_reg(131) <= "00000000001001110111000000000100";
         f_reg(132) <= "00000001111101011110000000000100";
         f_reg(133) <= "00010100110101000000000100100010";
         f_reg(134) <= "10101100000001100000010010100000";
         f_reg(135) <= "00000000000000000000000000000000";
         f_reg(136) <= "00000000000000000000000000000000";
         f_reg(137) <= "00000000000011000011100101000010";
         f_reg(138) <= "00000000000110101010100101000010";
         f_reg(139) <= "00010101100110100000000100011100";
         f_reg(140) <= "10101100000011000000010011011000";
         f_reg(141) <= "00000001110001100110000000100010";
         f_reg(142) <= "00000011100101001101000000100010";
         f_reg(143) <= "00000001011000110011000000100111";
         f_reg(144) <= "00000011001100011010000000100111";
         f_reg(145) <= "00010101101110110000000100010110";
         f_reg(146) <= "10101100000011010000010010100100";
         f_reg(147) <= "00000000011010010110100000100100";
         f_reg(148) <= "00000010001101111101100000100100";
         f_reg(149) <= "00000000100011100001100000100101";
         f_reg(150) <= "00000010010111001000100000100101";
         f_reg(151) <= "00000001000001110100100000100110";
         f_reg(152) <= "00000010110101011011100000100110";
         f_reg(153) <= "00111100000001000000101100011101";
         f_reg(154) <= "00111100000100100000101100011101";
         f_reg(155) <= "00000000100001110111000000100010";
         f_reg(156) <= "00000010010101011110000000100010";
         f_reg(157) <= "00000000000010000011100010000010";
         f_reg(158) <= "00000000000101101010100010000010";
         f_reg(159) <= "00000001110011100100000000000100";
         f_reg(160) <= "00000011100111001011000000000100";
         f_reg(161) <= "00010100110101000000000100000110";
         f_reg(162) <= "10101100000001100000010011011100";
         f_reg(163) <= "00000000000010000011000000100111";
         f_reg(164) <= "00000000000101101010000000100111";
         f_reg(165) <= "00010100110101000000000100000010";
         f_reg(166) <= "10101100000001100000010011100000";
         f_reg(167) <= "00101101001001101000101000001000";
         f_reg(168) <= "00101110111101001000101000001000";
         f_reg(169) <= "00000001101011000100100000100111";
         f_reg(170) <= "00000011011110101011100000100111";
         f_reg(171) <= "00010101100110100000000011111100";
         f_reg(172) <= "10101100000011000000010011100100";
         f_reg(173) <= "00000000111000100110000000100001";
         f_reg(174) <= "00000010101100001101000000100001";
         f_reg(175) <= "00111100000001110011100101100011";
         f_reg(176) <= "00111100000101010011100101100011";
         f_reg(177) <= "00000000110001000001000000100111";
         f_reg(178) <= "00000010100100101000000000100111";
         f_reg(179) <= "00010100010100000000000011110100";
         f_reg(180) <= "10101100000000100000010011101000";
         f_reg(181) <= "00000000000010100001001110000010";
         f_reg(182) <= "00000000000110001000001110000010";
         f_reg(183) <= "00000001101000000101000000100000";
         f_reg(184) <= "00000011011000001100000000100000";
         f_reg(185) <= "00000000000000000000000000000000";
         f_reg(186) <= "00000000000000000000000000000000";
         f_reg(187) <= "00100100100011011111100000101100";
         f_reg(188) <= "00100110010110111111100000101100";
         f_reg(189) <= "00101000110001000001110110011111";
         f_reg(190) <= "00101010100100100001110110011111";
         f_reg(191) <= "10001100000001100000010011011100";
         f_reg(192) <= "10001100000101000000010011011100";
         f_reg(193) <= "00010100110101001111111111111110";
         f_reg(194) <= "00010101000101100000000011100101";
         f_reg(195) <= "10101100000010000000010011011100";
         f_reg(196) <= "00000001110001100100000000100000";
         f_reg(197) <= "00000011100101001011000000100000";
         f_reg(198) <= "00000001011000110111000000100001";
         f_reg(199) <= "00000011001100011110000000100001";
         f_reg(200) <= "00000001101010000101100000100101";
         f_reg(201) <= "00000011011101101100100000100101";
         f_reg(202) <= "00000000010001110001100000000111";
         f_reg(203) <= "00000010000101011000100000000111";
         f_reg(204) <= "00000001001011000110100000100001";
         f_reg(205) <= "00000010111110101101100000100001";
         f_reg(206) <= "00000000000000000000000000000000";
         f_reg(207) <= "00000000000000000000000000000000";
         f_reg(208) <= "00101100001000010001100101111000";
         f_reg(209) <= "00101101111011110001100101111000";
         f_reg(210) <= "00010101010110000000000011010101";
         f_reg(211) <= "10101100000010100000010010101000";
         f_reg(212) <= "00000001011001010100000000100100";
         f_reg(213) <= "00000011001100111011000000100100";
         f_reg(214) <= "00010101000101100000000011010001";
         f_reg(215) <= "10101100000010000000010010101100";
         f_reg(216) <= "10001100000001110000010011011100";
         f_reg(217) <= "10001100000101010000010011011100";
         f_reg(218) <= "00010100111101011111111111111110";
         f_reg(219) <= "00000000111001000001000000100000";
         f_reg(220) <= "00000010101100101000000000100000";
         f_reg(221) <= "00000000010001100100100000100000";
         f_reg(222) <= "00000010000101001011100000100000";
         f_reg(223) <= "00000000000001100110011011000011";
         f_reg(224) <= "00000000000101001101011011000011";
         f_reg(225) <= "00000001110011000110000000000100";
         f_reg(226) <= "00000011100110101101000000000100";
         f_reg(227) <= "10001100000010100000010011100100";
         f_reg(228) <= "10001100000110000000010011100100";
         f_reg(229) <= "00010101010110001111111111111110";
         f_reg(230) <= "10001100000010110000010011011000";
         f_reg(231) <= "10001100000110010000010011011000";
         f_reg(232) <= "00010101011110011111111111111110";
         f_reg(233) <= "00000001010010110010100000101010";
         f_reg(234) <= "00000011000110011001100000101010";
         f_reg(235) <= "10001100000010000000010011100000";
         f_reg(236) <= "10001100000101100000010011100000";
         f_reg(237) <= "00010101000101101111111111111110";
         f_reg(238) <= "00000001000011010011100000101011";
         f_reg(239) <= "00000010110110111010100000101011";
         f_reg(240) <= "00010100110101000000000010110111";
         f_reg(241) <= "10101100000001100000010010110000";
         f_reg(242) <= "00110001100001001010010100111111";
         f_reg(243) <= "00110011010100101010010100111111";
         f_reg(244) <= "10001100000000100000010011101000";
         f_reg(245) <= "10001100000100000000010011101000";
         f_reg(246) <= "00010100010100001111111111111110";
         f_reg(247) <= "00000000011000100111000000000110";
         f_reg(248) <= "00000010001100001110000000000110";
         f_reg(249) <= "00000000111001010101000000100111";
         f_reg(250) <= "00000010101100111100000000100111";
         f_reg(251) <= "00100001010010111101011101010111";
         f_reg(252) <= "00100011000110011101011101010111";
         f_reg(253) <= "00101000100010000001110011001011";
         f_reg(254) <= "00101010010101100001110011001011";
         f_reg(255) <= "00010101110111000000000010101000";
         f_reg(256) <= "10101100000011100000010010110100";
         f_reg(257) <= "00010100101100110000000010100110";
         f_reg(258) <= "10101100000001010000010010111000";
         f_reg(259) <= "00010101001101110000000010100100";
         f_reg(260) <= "10101100000010010000010010111100";
         f_reg(261) <= "00010101110111000000000010100010";
         f_reg(262) <= "10101100000011100000010011000000";
         f_reg(263) <= "00111000111011011011111110101011";
         f_reg(264) <= "00111010101110111011111110101011";
         f_reg(265) <= "00101001011001101011000111001110";
         f_reg(266) <= "00101011001101001011000111001110";
         f_reg(267) <= "00010100001011110000000010011100";
         f_reg(268) <= "10101100000000010000010011000100";
         f_reg(269) <= "00010100110101000000000010011010";
         f_reg(270) <= "10101100000001100000010011001000";
         f_reg(271) <= "00100001101011000011010101111100";
         f_reg(272) <= "00100011011110100011010101111100";
         f_reg(273) <= "00010100011100010000000010010110";
         f_reg(274) <= "10101100000000110000010011001100";
         f_reg(275) <= "00000001100010110001000000100100";
         f_reg(276) <= "00000011010110011000000000100100";
         f_reg(277) <= "00100000010010100001001001100010";
         f_reg(278) <= "00100010000110000001001001100010";
         f_reg(279) <= "00010101000101100000000010010000";
         f_reg(280) <= "10101100000010000000010011010000";
         f_reg(281) <= "00010101010110000000000010001110";
         f_reg(282) <= "10101100000010100000010011010100";
         f_reg(283) <= "00100011110111011111111100000110";
         f_reg(284) <= "00010011101000000000000000100000";
         f_reg(285) <= "00100011110111011111111000001100";
         f_reg(286) <= "00010011101000000000000000011110";
         f_reg(287) <= "00100011110111011111110100010010";
         f_reg(288) <= "00010011101000000000000000011100";
         f_reg(289) <= "00100011110111101111111111111111";
         f_reg(290) <= "00100011111111111111111111111111";
         f_reg(291) <= "00010111110111110000000010000100";
         f_reg(292) <= "00011111111000001111111100110111";
         f_reg(293) <= "00010000000000000000000100001111";
         f_reg(294) <= "00000000000000000000000000000000";
         f_reg(295) <= "00000000000000000000000000000000";
         f_reg(296) <= "00000000000000000000000000000000";
         f_reg(297) <= "00000000000000000000000000000000";
         f_reg(298) <= "00000000000000000000000000000000";
         f_reg(299) <= "00000000000000000000000000000000";
         f_reg(300) <= "00000000000000000000000000000000";
         f_reg(301) <= "00000000000000000000000000000000";
         f_reg(302) <= "00000000000000000000000000000000";
         f_reg(303) <= "00000000000000000000000000000000";
         f_reg(304) <= "00000000000000000000000000000000";
         f_reg(305) <= "00000000000000000000000000000000";
         f_reg(306) <= "00000000000000000000000000000000";
         f_reg(307) <= "00000000000000000000000000000000";
         f_reg(308) <= "00000000000000000000000000000000";
         f_reg(309) <= "00000000000000000000000000000000";
         f_reg(310) <= "00000000000000000000000000000000";
         f_reg(311) <= "00000000000000000000000000000000";
         f_reg(312) <= "00000000000000000000000000000000";
         f_reg(313) <= "00000000000000000000000000000000";
         f_reg(314) <= "00000000000000000000000000000000";
         f_reg(315) <= "00000000000000000000000000000000";
         f_reg(316) <= "10001100000111010000100001000000";
         f_reg(317) <= "00011111101000000000000000000011";
         f_reg(318) <= "00100000000111010000000000111100";
         f_reg(319) <= "00010000000000000000000000000010";
         f_reg(320) <= "00100000000111010000000000000000";
         f_reg(321) <= "00010100001011110000000001100110";
         f_reg(322) <= "10101111101000010000011111001000";
         f_reg(323) <= "10001100000111010000100001000000";
         f_reg(324) <= "00011111101000000000000000000011";
         f_reg(325) <= "00100000000111010000000000111100";
         f_reg(326) <= "00010000000000000000000000000010";
         f_reg(327) <= "00100000000111010000000000000000";
         f_reg(328) <= "00010100010100000000000001011111";
         f_reg(329) <= "10101111101000100000011111001100";
         f_reg(330) <= "10001100000111010000100001000000";
         f_reg(331) <= "00011111101000000000000000000011";
         f_reg(332) <= "00100000000111010000000000111100";
         f_reg(333) <= "00010000000000000000000000000010";
         f_reg(334) <= "00100000000111010000000000000000";
         f_reg(335) <= "00010100011100010000000001011000";
         f_reg(336) <= "10101111101000110000011111010000";
         f_reg(337) <= "10001100000111010000100001000000";
         f_reg(338) <= "00011111101000000000000000000011";
         f_reg(339) <= "00100000000111010000000000111100";
         f_reg(340) <= "00010000000000000000000000000010";
         f_reg(341) <= "00100000000111010000000000000000";
         f_reg(342) <= "00010100100100100000000001010001";
         f_reg(343) <= "10101111101001000000011111010100";
         f_reg(344) <= "10001100000111010000100001000000";
         f_reg(345) <= "00011111101000000000000000000011";
         f_reg(346) <= "00100000000111010000000000111100";
         f_reg(347) <= "00010000000000000000000000000010";
         f_reg(348) <= "00100000000111010000000000000000";
         f_reg(349) <= "00010100101100110000000001001010";
         f_reg(350) <= "10101111101001010000011111011000";
         f_reg(351) <= "10001100000111010000100001000000";
         f_reg(352) <= "00011111101000000000000000000011";
         f_reg(353) <= "00100000000111010000000000111100";
         f_reg(354) <= "00010000000000000000000000000010";
         f_reg(355) <= "00100000000111010000000000000000";
         f_reg(356) <= "00010100110101000000000001000011";
         f_reg(357) <= "10101111101001100000011111011100";
         f_reg(358) <= "10001100000111010000100001000000";
         f_reg(359) <= "00011111101000000000000000000011";
         f_reg(360) <= "00100000000111010000000000111100";
         f_reg(361) <= "00010000000000000000000000000010";
         f_reg(362) <= "00100000000111010000000000000000";
         f_reg(363) <= "00010100111101010000000000111100";
         f_reg(364) <= "10101111101001110000011111100000";
         f_reg(365) <= "10001100000111010000100001000000";
         f_reg(366) <= "00011111101000000000000000000011";
         f_reg(367) <= "00100000000111010000000000111100";
         f_reg(368) <= "00010000000000000000000000000010";
         f_reg(369) <= "00100000000111010000000000000000";
         f_reg(370) <= "00010101000101100000000000110101";
         f_reg(371) <= "10101111101010000000011111100100";
         f_reg(372) <= "10001100000111010000100001000000";
         f_reg(373) <= "00011111101000000000000000000011";
         f_reg(374) <= "00100000000111010000000000111100";
         f_reg(375) <= "00010000000000000000000000000010";
         f_reg(376) <= "00100000000111010000000000000000";
         f_reg(377) <= "00010101001101110000000000101110";
         f_reg(378) <= "10101111101010010000011111101000";
         f_reg(379) <= "10001100000111010000100001000000";
         f_reg(380) <= "00011111101000000000000000000011";
         f_reg(381) <= "00100000000111010000000000111100";
         f_reg(382) <= "00010000000000000000000000000010";
         f_reg(383) <= "00100000000111010000000000000000";
         f_reg(384) <= "00010101010110000000000000100111";
         f_reg(385) <= "10101111101010100000011111101100";
         f_reg(386) <= "10001100000111010000100001000000";
         f_reg(387) <= "00011111101000000000000000000011";
         f_reg(388) <= "00100000000111010000000000111100";
         f_reg(389) <= "00010000000000000000000000000010";
         f_reg(390) <= "00100000000111010000000000000000";
         f_reg(391) <= "00010101011110010000000000100000";
         f_reg(392) <= "10101111101010110000011111110000";
         f_reg(393) <= "10001100000111010000100001000000";
         f_reg(394) <= "00011111101000000000000000000011";
         f_reg(395) <= "00100000000111010000000000111100";
         f_reg(396) <= "00010000000000000000000000000010";
         f_reg(397) <= "00100000000111010000000000000000";
         f_reg(398) <= "00010101100110100000000000011001";
         f_reg(399) <= "10101111101011000000011111110100";
         f_reg(400) <= "10001100000111010000100001000000";
         f_reg(401) <= "00011111101000000000000000000011";
         f_reg(402) <= "00100000000111010000000000111100";
         f_reg(403) <= "00010000000000000000000000000010";
         f_reg(404) <= "00100000000111010000000000000000";
         f_reg(405) <= "00010101101110110000000000010010";
         f_reg(406) <= "10101111101011010000011111111000";
         f_reg(407) <= "10001100000111010000100001000000";
         f_reg(408) <= "00011111101000000000000000000011";
         f_reg(409) <= "00100000000111010000000000111100";
         f_reg(410) <= "00010000000000000000000000000010";
         f_reg(411) <= "00100000000111010000000000000000";
         f_reg(412) <= "00010101110111000000000000001011";
         f_reg(413) <= "10101111101011100000011111111100";
         f_reg(414) <= "10001100000111010000100001000000";
         f_reg(415) <= "00011111101000000000000000000011";
         f_reg(416) <= "00100000000111010000000000111100";
         f_reg(417) <= "00010000000000000000000000000010";
         f_reg(418) <= "00100000000111010000000000000000";
         f_reg(419) <= "00010111110111110000000000000100";
         f_reg(420) <= "10101111101111100000100000000000";
         f_reg(421) <= "10101100000111010000100001000000";
         f_reg(422) <= "00010000000000001111111101111011";
         f_reg(423) <= "10001100000111010000100001000000";
         f_reg(424) <= "10001111101000010000011111001000";
         f_reg(425) <= "10001100000111010000100001000000";
         f_reg(426) <= "10001111101011110000011111001000";
         f_reg(427) <= "00010100001011111111111111111100";
         f_reg(428) <= "10001100000111010000100001000000";
         f_reg(429) <= "10001111101000100000011111001100";
         f_reg(430) <= "10001100000111010000100001000000";
         f_reg(431) <= "10001111101100000000011111001100";
         f_reg(432) <= "00010100010100001111111111111100";
         f_reg(433) <= "10001100000111010000100001000000";
         f_reg(434) <= "10001111101000110000011111010000";
         f_reg(435) <= "10001100000111010000100001000000";
         f_reg(436) <= "10001111101100010000011111010000";
         f_reg(437) <= "00010100011100011111111111111100";
         f_reg(438) <= "10001100000111010000100001000000";
         f_reg(439) <= "10001111101001000000011111010100";
         f_reg(440) <= "10001100000111010000100001000000";
         f_reg(441) <= "10001111101100100000011111010100";
         f_reg(442) <= "00010100100100101111111111111100";
         f_reg(443) <= "10001100000111010000100001000000";
         f_reg(444) <= "10001111101001010000011111011000";
         f_reg(445) <= "10001100000111010000100001000000";
         f_reg(446) <= "10001111101100110000011111011000";
         f_reg(447) <= "00010100101100111111111111111100";
         f_reg(448) <= "10001100000111010000100001000000";
         f_reg(449) <= "10001111101001100000011111011100";
         f_reg(450) <= "10001100000111010000100001000000";
         f_reg(451) <= "10001111101101000000011111011100";
         f_reg(452) <= "00010100110101001111111111111100";
         f_reg(453) <= "10001100000111010000100001000000";
         f_reg(454) <= "10001111101001110000011111100000";
         f_reg(455) <= "10001100000111010000100001000000";
         f_reg(456) <= "10001111101101010000011111100000";
         f_reg(457) <= "00010100111101011111111111111100";
         f_reg(458) <= "10001100000111010000100001000000";
         f_reg(459) <= "10001111101010000000011111100100";
         f_reg(460) <= "10001100000111010000100001000000";
         f_reg(461) <= "10001111101101100000011111100100";
         f_reg(462) <= "00010101000101101111111111111100";
         f_reg(463) <= "10001100000111010000100001000000";
         f_reg(464) <= "10001111101010010000011111101000";
         f_reg(465) <= "10001100000111010000100001000000";
         f_reg(466) <= "10001111101101110000011111101000";
         f_reg(467) <= "00010101001101111111111111111100";
         f_reg(468) <= "10001100000111010000100001000000";
         f_reg(469) <= "10001111101010100000011111101100";
         f_reg(470) <= "10001100000111010000100001000000";
         f_reg(471) <= "10001111101110000000011111101100";
         f_reg(472) <= "00010101010110001111111111111100";
         f_reg(473) <= "10001100000111010000100001000000";
         f_reg(474) <= "10001111101010110000011111110000";
         f_reg(475) <= "10001100000111010000100001000000";
         f_reg(476) <= "10001111101110010000011111110000";
         f_reg(477) <= "00010101011110011111111111111100";
         f_reg(478) <= "10001100000111010000100001000000";
         f_reg(479) <= "10001111101011000000011111110100";
         f_reg(480) <= "10001100000111010000100001000000";
         f_reg(481) <= "10001111101110100000011111110100";
         f_reg(482) <= "00010101100110101111111111111100";
         f_reg(483) <= "10001100000111010000100001000000";
         f_reg(484) <= "10001111101011010000011111111000";
         f_reg(485) <= "10001100000111010000100001000000";
         f_reg(486) <= "10001111101110110000011111111000";
         f_reg(487) <= "00010101101110111111111111111100";
         f_reg(488) <= "10001100000111010000100001000000";
         f_reg(489) <= "10001111101011100000011111111100";
         f_reg(490) <= "10001100000111010000100001000000";
         f_reg(491) <= "10001111101111000000011111111100";
         f_reg(492) <= "00010101110111001111111111111100";
         f_reg(493) <= "10001100000111010000100001000000";
         f_reg(494) <= "10001111101111100000100000000000";
         f_reg(495) <= "10001100000111010000100001000000";
         f_reg(496) <= "10001111101111110000100000000000";
         f_reg(497) <= "00010111110111111111111111111100";
         f_reg(498) <= "00010000000000001111111100101111";
         f_reg(499) <= "00000000000000000000000000000000";
         f_reg(500) <= "00000000000000000000000000000000";
         f_reg(501) <= "00000000000000000000000000000000";
         f_reg(502) <= "00000000000000000000000000000000";
         f_reg(503) <= "00000000000000000000000000000000";
         f_reg(504) <= "00000000000000000000000000000000";
         f_reg(505) <= "00000000000000000000000000000000";
         f_reg(506) <= "00000000000000000000000000000000";
         f_reg(507) <= "00000000000000000000000000000000";
         f_reg(508) <= "00000000000000000000000000000000";
         f_reg(509) <= "00000000000000000000000000000000";
         f_reg(510) <= "00000000000000000000000000000000";
         f_reg(511) <= "00000000000000000000000000000000";
         f_reg(512) <= "00000000000000000000000000000000";
         f_reg(513) <= "00000000000000000000000000000000";
         f_reg(514) <= "00000000000000000000000000000000";
         f_reg(515) <= "00000000000000000000000000000000";
         f_reg(516) <= "00000000000000000000000000000000";
         f_reg(517) <= "00000000000000000000000000000000";
         f_reg(518) <= "00000000000000000000000000000000";
         f_reg(519) <= "00000000000000000000000000000000";
         f_reg(520) <= "00000000000000000000000000000000";
         f_reg(521) <= "00000000000000000000000000000000";
         f_reg(522) <= "00000000000000000000000000000000";
         f_reg(523) <= "00000000000000000000000000000000";
         f_reg(524) <= "00000000000000000000000000000000";
         f_reg(525) <= "00000000000000000000000000000000";
         f_reg(526) <= "00000000000000000000000000000000";
         f_reg(527) <= "00000000000000000000000000000000";
         f_reg(528) <= "00000000000000000000000000000000";
         f_reg(529) <= "00000000000000000000001111100111";
         f_reg(530) <= "00000000000000000000000000000000";
         f_reg(531) <= "00000000000000000000000000000000";
         f_reg(532) <= "00000000000000000000000000000000";
         f_reg(533) <= "00000000000000000000000000000000";
         f_reg(534) <= "00000000000000000000000000000000";
         f_reg(535) <= "00000000000000000000000000000000";
         f_reg(536) <= "00000000000000000000000000000000";
         f_reg(537) <= "00000000000000000000000000000000";
         f_reg(538) <= "00000000000000000000000000000000";
         f_reg(539) <= "00000000000000000000000000000000";
         f_reg(540) <= "00000000000000000000000000000000";
         f_reg(541) <= "00000000000000000000000000000000";
         f_reg(542) <= "00000000000000000000000000000000";
         f_reg(543) <= "00000000000000000000000000000000";
         f_reg(544) <= "00000000000000000000000000000000";
         f_reg(545) <= "00000000000000000000000000000000";
         f_reg(546) <= "00000000000000000000000000000000";
         f_reg(547) <= "00000000000000000000000000000000";
         f_reg(548) <= "00000000000000000000000000000000";
         f_reg(549) <= "00000000000000000000000000000000";
         f_reg(550) <= "00000000000000000000000000000000";
         f_reg(551) <= "00000000000000000000000000000000";
         f_reg(552) <= "00000000000000000000000000000000";
         f_reg(553) <= "00000000000000000000000000000000";
         f_reg(554) <= "00000000000000000000000000000000";
         f_reg(555) <= "00000000000000000000000000000000";
         f_reg(556) <= "00000000000000000000000000000000";
         f_reg(557) <= "00000000000000000000000000000000";
         f_reg(558) <= "00000000000000000000000000000000";
         f_reg(559) <= "00000000000000000000000000000000";
         f_reg(560) <= "00000000000000000000000000000000";
         f_reg(561) <= "00000000000000000000000000000000";
         f_reg(562) <= "00000000000000000000000000000000";
         f_reg(563) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 3914
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- XORI R2 R0 -13506
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- SW R1 R0 1172
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SRL R3 R0 20
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SUBU R4 R1 R2
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- XORI R5 R2 11459
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- ANDI R6 R4 23545
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- ADD R7 R2 R6
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- SUB R8 R3 R2
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- ADDIU R9 R4 -9117
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- ANDI R10 R3 7716
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- SRLV R11 R8 R8
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- SW R6 R0 1176
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- ADD R12 R6 R9
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- ADD R13 R9 R8
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- SRLV R14 R12 R1
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SRLV R15 R10 R14
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- SLTI R16 R11 11687
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- SW R1 R0 1180
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- SRLV R17 R4 R9
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- SLLV R18 R7 R1
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- SW R6 R0 1184
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- NOP
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- SRL R19 R12 5
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- SUB R20 R18 R6
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- NOR R21 R11 R16
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- SW R13 R0 1188
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- AND R22 R16 R9
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- OR R23 R4 R18
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- XOR R24 R17 R19
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- LUI R25 2845
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- SUB R26 R25 R19
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- SRL R27 R17 2
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- SLLV R28 R26 R26
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- NOR R29 R0 R28
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- SLTIU R30 R24 -30200
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- NOR R2 R22 R20
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- ADDU R3 R27 R15
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- LUI R8 14691
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- NOR R14 R30 R25
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SRL R7 R10 14
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- ADD R6 R22 R0
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- NOP
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- ADDIU R13 R25 -2004
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- SLTI R16 R30 7583
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- ADD R9 R26 R21
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- ADDU R4 R11 R23
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- OR R18 R13 R9
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- SRAV R19 R8 R7
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- ADDU R17 R2 R3
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- NOP
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SLTIU R1 R1 6520
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SW R6 R0 1192
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- AND R24 R18 R5
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SW R24 R0 1196
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- ADD R27 R28 R16
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- ADD R15 R27 R21
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- SRA R10 R21 27
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- SLLV R10 R10 R4
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- SLT R22 R20 R12
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- SLTU R25 R29 R17
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- SW R21 R0 1200
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- ANDI R30 R10 -23233
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- SRLV R26 R14 R19
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- NOR R11 R25 R22
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- ADDI R23 R11 -10409
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- SLTI R13 R30 7371
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SW R26 R0 1204
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- SW R22 R0 1208
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- SW R15 R0 1212
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SW R26 R0 1216
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- XORI R9 R25 -16469
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- SLTI R8 R23 -20018
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- SW R1 R0 1220
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- SW R8 R0 1224
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- ADDI R7 R9 13692
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- SW R19 R0 1228
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- AND R2 R7 R23
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- ADDI R3 R2 4706
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- SW R13 R0 1232
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SW R3 R0 1236
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- BGTZ R31 -82
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- BEQ R0 R0 478
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- LUI R30 999
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- LUI R31 999
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- LUI R1 3914
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- LUI R15 3914
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- XORI R2 R0 -13506
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- XORI R16 R0 -13506
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- BNE R1 R15 328
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- SW R1 R0 1172
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SRL R3 R0 20
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SRL R17 R0 20
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- SUBU R4 R1 R2
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- SUBU R18 R15 R16
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- XORI R5 R2 11459
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- XORI R19 R16 11459
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- ANDI R6 R4 23545
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- ANDI R20 R18 23545
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- ADD R7 R2 R6
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- ADD R21 R16 R20
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- SUB R8 R3 R2
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- SUB R22 R17 R16
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- ADDIU R9 R4 -9117
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- ADDIU R23 R18 -9117
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- ANDI R10 R3 7716
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- ANDI R24 R17 7716
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- SRLV R11 R8 R8
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- SRLV R25 R22 R22
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- BNE R6 R20 308
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- SW R6 R0 1176
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- ADD R12 R6 R9
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- ADD R26 R20 R23
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- ADD R13 R9 R8
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- ADD R27 R23 R22
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- SRLV R14 R12 R1
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- SRLV R28 R26 R15
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- SRLV R2 R10 R14
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SRLV R16 R24 R28
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- SLTI R3 R11 11687
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- SLTI R17 R25 11687
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- BNE R1 R15 296
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SW R1 R0 1180
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- SRLV R8 R4 R9
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- SRLV R22 R18 R23
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- SLLV R14 R7 R1
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- SLLV R28 R21 R15
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- BNE R6 R20 290
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- SW R6 R0 1184
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- NOP
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- NOP
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- SRL R7 R12 5
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SRL R21 R26 5
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- BNE R12 R26 284
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- SW R12 R0 1240
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- SUB R12 R14 R6
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- SUB R26 R28 R20
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- NOR R6 R11 R3
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- NOR R20 R25 R17
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- BNE R13 R27 278
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- SW R13 R0 1188
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- AND R13 R3 R9
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- AND R27 R17 R23
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- OR R3 R4 R14
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- OR R17 R18 R28
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- XOR R9 R8 R7
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- XOR R23 R22 R21
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- LUI R4 2845
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- LUI R18 2845
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- SUB R14 R4 R7
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- SUB R28 R18 R21
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- SRL R7 R8 2
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- SRL R21 R22 2
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- SLLV R8 R14 R14
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- SLLV R22 R28 R28
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- BNE R6 R20 262
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- SW R6 R0 1244
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- NOR R6 R0 R8
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- NOR R20 R0 R22
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- BNE R6 R20 258
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- SW R6 R0 1248
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- SLTIU R6 R9 -30200
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- SLTIU R20 R23 -30200
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- NOR R9 R13 R12
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- NOR R23 R27 R26
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- BNE R12 R26 252
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- SW R12 R0 1252
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- ADDU R12 R7 R2
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- ADDU R26 R21 R16
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- LUI R7 14691
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- LUI R21 14691
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- NOR R2 R6 R4
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- NOR R16 R20 R18
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- BNE R2 R16 244
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- SW R2 R0 1256
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- SRL R2 R10 14
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SRL R16 R24 14
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- ADD R10 R13 R0
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- ADD R24 R27 R0
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- NOP
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- NOP
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- ADDIU R13 R4 -2004
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- ADDIU R27 R18 -2004
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- SLTI R4 R6 7583
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- SLTI R18 R20 7583
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- LW R6 R0 1244
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- LW R20 R0 1244
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- BNE R6 R20 -2
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- BNE R8 R22 229
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- SW R8 R0 1244
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- ADD R8 R14 R6
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- ADD R22 R28 R20
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- ADDU R14 R11 R3
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- ADDU R28 R25 R17
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- OR R11 R13 R8
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- OR R25 R27 R22
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- SRAV R3 R7 R2
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- SRAV R17 R21 R16
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- ADDU R13 R9 R12
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- ADDU R27 R23 R26
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- NOP
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- NOP
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- SLTIU R1 R1 6520
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- SLTIU R15 R15 6520
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- BNE R10 R24 213
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- SW R10 R0 1192
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- AND R8 R11 R5
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- AND R22 R25 R19
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- BNE R8 R22 209
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- SW R8 R0 1196
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- LW R7 R0 1244
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- LW R21 R0 1244
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- BNE R7 R21 -2
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- ADD R2 R7 R4
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- ADD R16 R21 R18
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- ADD R9 R2 R6
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- ADD R23 R16 R20
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- SRA R12 R6 27
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- SRA R26 R20 27
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- SLLV R12 R12 R14
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- SLLV R26 R26 R28
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- LW R10 R0 1252
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- LW R24 R0 1252
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- BNE R10 R24 -2
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- LW R11 R0 1240
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- LW R25 R0 1240
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- BNE R11 R25 -2
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- SLT R5 R10 R11
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- SLT R19 R24 R25
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- LW R8 R0 1248
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- LW R22 R0 1248
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- BNE R8 R22 -2
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- SLTU R7 R8 R13
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- SLTU R21 R22 R27
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- BNE R6 R20 183
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- SW R6 R0 1200
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- ANDI R4 R12 -23233
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- ANDI R18 R26 -23233
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- LW R2 R0 1256
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- LW R16 R0 1256
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- BNE R2 R16 -2
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- SRLV R14 R2 R3
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- SRLV R28 R16 R17
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- NOR R10 R7 R5
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- NOR R24 R21 R19
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- ADDI R11 R10 -10409
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- ADDI R25 R24 -10409
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- SLTI R8 R4 7371
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- SLTI R22 R18 7371
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- BNE R14 R28 168
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- SW R14 R0 1204
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- BNE R5 R19 166
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- SW R5 R0 1208
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- BNE R9 R23 164
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- SW R9 R0 1212
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- BNE R14 R28 162
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- SW R14 R0 1216
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- XORI R13 R7 -16469
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- XORI R27 R21 -16469
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- SLTI R6 R11 -20018
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- SLTI R20 R25 -20018
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- BNE R1 R15 156
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- SW R1 R0 1220
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- BNE R6 R20 154
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- SW R6 R0 1224
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- ADDI R12 R13 13692
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- ADDI R26 R27 13692
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- BNE R3 R17 150
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- SW R3 R0 1228
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- AND R2 R12 R11
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- AND R16 R26 R25
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- ADDI R10 R2 4706
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- ADDI R24 R16 4706
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- BNE R8 R22 144
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- SW R8 R0 1232
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- BNE R10 R24 142
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- SW R10 R0 1236
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- BEQ R29 R0 32
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- BEQ R29 R0 30
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- BEQ R29 R0 28
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- BNE R30 R31 132
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- BGTZ R31 -201
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- BEQ R0 R0 271
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- NOP
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- NOP
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- NOP
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- NOP
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- NOP
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- NOP
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- NOP
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- NOP
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- NOP
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- NOP
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- NOP
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- NOP
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- NOP
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- NOP
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- NOP
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- NOP
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- NOP
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- NOP
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- NOP
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- NOP
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- NOP
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- NOP
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- SW R1 R29 1992
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- SW R2 R29 1996
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- SW R3 R29 2000
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- SW R4 R29 2004
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- SW R5 R29 2008
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- SW R6 R29 2012
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- SW R7 R29 2016
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- SW R8 R29 2020
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- SW R9 R29 2024
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- SW R10 R29 2028
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- SW R11 R29 2032
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- SW R12 R29 2036
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- SW R13 R29 2040
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- SW R14 R29 2044
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- SW R30 R29 2048
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- SW R29 R0 2112
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- BEQ R0 R0 -133
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- LW R1 R29 1992
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R15 R29 1992
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- LW R2 R29 1996
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- LW R16 R29 1996
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- LW R3 R29 2000
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- LW R17 R29 2000
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- LW R4 R29 2004
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- LW R18 R29 2004
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- LW R5 R29 2008
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- LW R19 R29 2008
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- LW R6 R29 2012
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- LW R20 R29 2012
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- LW R7 R29 2016
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- LW R21 R29 2016
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- LW R8 R29 2020
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- LW R22 R29 2020
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- LW R9 R29 2024
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- LW R23 R29 2024
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- LW R10 R29 2028
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- LW R24 R29 2028
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- LW R11 R29 2032
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- LW R25 R29 2032
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- LW R12 R29 2036
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- LW R26 R29 2036
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- LW R13 R29 2040
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- LW R27 R29 2040
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- LW R14 R29 2044
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- LW R28 R29 2044
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- LW R30 R29 2048
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- LW R29 R0 2112
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- LW R31 R29 2048
                        f_data <= f_reg(496);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(497) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(497);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(498) =>
                        -- BEQ R0 R0 -209
                        f_data <= f_reg(498);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(499) =>
                        -- NOP
                        f_data <= f_reg(499);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(500) =>
                        -- NOP
                        f_data <= f_reg(500);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(501) =>
                        -- NOP
                        f_data <= f_reg(501);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(502) =>
                        -- NOP
                        f_data <= f_reg(502);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(503) =>
                        -- NOP
                        f_data <= f_reg(503);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(504) =>
                        -- NOP
                        f_data <= f_reg(504);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(505) =>
                        -- NOP
                        f_data <= f_reg(505);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(506) =>
                        -- NOP
                        f_data <= f_reg(506);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(507) =>
                        -- NOP
                        f_data <= f_reg(507);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(508) =>
                        -- NOP
                        f_data <= f_reg(508);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(509) =>
                        -- NOP
                        f_data <= f_reg(509);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(510) =>
                        -- NOP
                        f_data <= f_reg(510);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(511) =>
                        -- NOP
                        f_data <= f_reg(511);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(512) =>
                        -- NOP
                        f_data <= f_reg(512);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(513) =>
                        -- NOP
                        f_data <= f_reg(513);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(514) =>
                        -- NOP
                        f_data <= f_reg(514);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(515) =>
                        -- NOP
                        f_data <= f_reg(515);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(516) =>
                        -- NOP
                        f_data <= f_reg(516);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(517) =>
                        -- NOP
                        f_data <= f_reg(517);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(518) =>
                        -- NOP
                        f_data <= f_reg(518);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(519) =>
                        -- NOP
                        f_data <= f_reg(519);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(520) =>
                        -- NOP
                        f_data <= f_reg(520);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(521) =>
                        -- NOP
                        f_data <= f_reg(521);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(522) =>
                        -- NOP
                        f_data <= f_reg(522);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(523) =>
                        -- NOP
                        f_data <= f_reg(523);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(524) =>
                        -- NOP
                        f_data <= f_reg(524);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(525) =>
                        -- NOP
                        f_data <= f_reg(525);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(526) =>
                        -- NOP
                        f_data <= f_reg(526);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(527) =>
                        -- NOP
                        f_data <= f_reg(527);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(528) =>
                        -- NOP
                        f_data <= f_reg(528);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(529) =>
                        -- NOP
                        f_data <= f_reg(529);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(530) =>
                        -- NOP
                        f_data <= f_reg(530);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(531) =>
                        -- NOP
                        f_data <= f_reg(531);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(532) =>
                        -- NOP
                        f_data <= f_reg(532);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(533) =>
                        -- NOP
                        f_data <= f_reg(533);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(534) =>
                        -- NOP
                        f_data <= f_reg(534);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(535) =>
                        -- NOP
                        f_data <= f_reg(535);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(536) =>
                        -- NOP
                        f_data <= f_reg(536);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(537) =>
                        -- NOP
                        f_data <= f_reg(537);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(538) =>
                        -- NOP
                        f_data <= f_reg(538);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(539) =>
                        -- NOP
                        f_data <= f_reg(539);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(540) =>
                        -- NOP
                        f_data <= f_reg(540);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(541) =>
                        -- NOP
                        f_data <= f_reg(541);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(542) =>
                        -- NOP
                        f_data <= f_reg(542);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(543) =>
                        -- NOP
                        f_data <= f_reg(543);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(544) =>
                        -- NOP
                        f_data <= f_reg(544);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(545) =>
                        -- NOP
                        f_data <= f_reg(545);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(546) =>
                        -- NOP
                        f_data <= f_reg(546);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(547) =>
                        -- NOP
                        f_data <= f_reg(547);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(548) =>
                        -- NOP
                        f_data <= f_reg(548);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(549) =>
                        -- NOP
                        f_data <= f_reg(549);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(550) =>
                        -- NOP
                        f_data <= f_reg(550);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(551) =>
                        -- NOP
                        f_data <= f_reg(551);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(552) =>
                        -- NOP
                        f_data <= f_reg(552);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(553) =>
                        -- NOP
                        f_data <= f_reg(553);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(554) =>
                        -- NOP
                        f_data <= f_reg(554);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(555) =>
                        -- NOP
                        f_data <= f_reg(555);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(556) =>
                        -- NOP
                        f_data <= f_reg(556);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(557) =>
                        -- NOP
                        f_data <= f_reg(557);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(558) =>
                        -- NOP
                        f_data <= f_reg(558);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(559) =>
                        -- NOP
                        f_data <= f_reg(559);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(560) =>
                        -- NOP
                        f_data <= f_reg(560);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(561) =>
                        -- NOP
                        f_data <= f_reg(561);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(562) =>
                        -- NOP
                        f_data <= f_reg(562);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(563) =>
                        -- NOP
                        f_data <= f_reg(563);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(564) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010000111101001010";
                        f_reg(4) <= "00111000000000101100101100111110";
                        f_reg(5) <= "10101100000000010000010010010100";
                        f_reg(6) <= "00000000000000000001110100000010";
                        f_reg(7) <= "00000000001000100010000000100011";
                        f_reg(8) <= "00111000010001010010110011000011";
                        f_reg(9) <= "00110000100001100101101111111001";
                        f_reg(10) <= "00000000010001100011100000100000";
                        f_reg(11) <= "00000000011000100100000000100010";
                        f_reg(12) <= "00100100100010011101110001100011";
                        f_reg(13) <= "00110000011010100001111000100100";
                        f_reg(14) <= "00000001000010000101100000000110";
                        f_reg(15) <= "10101100000001100000010010011000";
                        f_reg(16) <= "00000000110010010110000000100000";
                        f_reg(17) <= "00000001001010000110100000100000";
                        f_reg(18) <= "00000000001011000111000000000110";
                        f_reg(19) <= "00000001110010100111100000000110";
                        f_reg(20) <= "00101001011100000010110110100111";
                        f_reg(21) <= "10101100000000010000010010011100";
                        f_reg(22) <= "00000001001001001000100000000110";
                        f_reg(23) <= "00000000001001111001000000000100";
                        f_reg(24) <= "10101100000001100000010010100000";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00000000000011001001100101000010";
                        f_reg(27) <= "00000010010001101010000000100010";
                        f_reg(28) <= "00000001011100001010100000100111";
                        f_reg(29) <= "10101100000011010000010010100100";
                        f_reg(30) <= "00000010000010011011000000100100";
                        f_reg(31) <= "00000000100100101011100000100101";
                        f_reg(32) <= "00000010001100111100000000100110";
                        f_reg(33) <= "00111100000110010000101100011101";
                        f_reg(34) <= "00000011001100111101000000100010";
                        f_reg(35) <= "00000000000100011101100010000010";
                        f_reg(36) <= "00000011010110101110000000000100";
                        f_reg(37) <= "00000000000111001110100000100111";
                        f_reg(38) <= "00101111000111101000101000001000";
                        f_reg(39) <= "00000010110101000001000000100111";
                        f_reg(40) <= "00000011011011110001100000100001";
                        f_reg(41) <= "00111100000010000011100101100011";
                        f_reg(42) <= "00000011110110010111000000100111";
                        f_reg(43) <= "00000000000010100011101110000010";
                        f_reg(44) <= "00000010110000000011000000100000";
                        f_reg(45) <= "00000000000000000000000000000000";
                        f_reg(46) <= "00100111001011011111100000101100";
                        f_reg(47) <= "00101011110100000001110110011111";
                        f_reg(48) <= "00000011010101010100100000100000";
                        f_reg(49) <= "00000001011101110010000000100001";
                        f_reg(50) <= "00000001101010011001000000100101";
                        f_reg(51) <= "00000000111010001001100000000111";
                        f_reg(52) <= "00000000010000111000100000100001";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00101100001000010001100101111000";
                        f_reg(55) <= "10101100000001100000010010101000";
                        f_reg(56) <= "00000010010001011100000000100100";
                        f_reg(57) <= "10101100000110000000010010101100";
                        f_reg(58) <= "00000011100100001101100000100000";
                        f_reg(59) <= "00000011011101010111100000100000";
                        f_reg(60) <= "00000000000101010101011011000011";
                        f_reg(61) <= "00000000100010100101000000000100";
                        f_reg(62) <= "00000010100011001011000000101010";
                        f_reg(63) <= "00000011101100011100100000101011";
                        f_reg(64) <= "10101100000101010000010010110000";
                        f_reg(65) <= "00110001010111101010010100111111";
                        f_reg(66) <= "00000010011011101101000000000110";
                        f_reg(67) <= "00000011001101100101100000100111";
                        f_reg(68) <= "00100001011101111101011101010111";
                        f_reg(69) <= "00101011110011010001110011001011";
                        f_reg(70) <= "10101100000110100000010010110100";
                        f_reg(71) <= "10101100000101100000010010111000";
                        f_reg(72) <= "10101100000011110000010010111100";
                        f_reg(73) <= "10101100000110100000010011000000";
                        f_reg(74) <= "00111011001010011011111110101011";
                        f_reg(75) <= "00101010111010001011000111001110";
                        f_reg(76) <= "10101100000000010000010011000100";
                        f_reg(77) <= "10101100000010000000010011001000";
                        f_reg(78) <= "00100001001001110011010101111100";
                        f_reg(79) <= "10101100000100110000010011001100";
                        f_reg(80) <= "00000000111101110001000000100100";
                        f_reg(81) <= "00100000010000110001001001100010";
                        f_reg(82) <= "10101100000011010000010011010000";
                        f_reg(83) <= "10101100000000110000010011010100";
                        f_reg(84) <= "00100011111111111111111111111111";
                        f_reg(85) <= "00011111111000001111111110101110";
                        f_reg(86) <= "00010000000000000000000111011110";
                        f_reg(87) <= "00111100000111100000001111100111";
                        f_reg(88) <= "00111100000111110000001111100111";
                        f_reg(89) <= "00000000000111101111010000000010";
                        f_reg(90) <= "00000000000111111111110000000010";
                        f_reg(91) <= "00111100000000010000111101001010";
                        f_reg(92) <= "00111100000011110000111101001010";
                        f_reg(93) <= "00111000000000101100101100111110";
                        f_reg(94) <= "00111000000100001100101100111110";
                        f_reg(95) <= "00010100001011110000000101001000";
                        f_reg(96) <= "10101100000000010000010010010100";
                        f_reg(97) <= "00000000000000000001110100000010";
                        f_reg(98) <= "00000000000000001000110100000010";
                        f_reg(99) <= "00000000001000100010000000100011";
                        f_reg(100) <= "00000001111100001001000000100011";
                        f_reg(101) <= "00111000010001010010110011000011";
                        f_reg(102) <= "00111010000100110010110011000011";
                        f_reg(103) <= "00110000100001100101101111111001";
                        f_reg(104) <= "00110010010101000101101111111001";
                        f_reg(105) <= "00000000010001100011100000100000";
                        f_reg(106) <= "00000010000101001010100000100000";
                        f_reg(107) <= "00000000011000100100000000100010";
                        f_reg(108) <= "00000010001100001011000000100010";
                        f_reg(109) <= "00100100100010011101110001100011";
                        f_reg(110) <= "00100110010101111101110001100011";
                        f_reg(111) <= "00110000011010100001111000100100";
                        f_reg(112) <= "00110010001110000001111000100100";
                        f_reg(113) <= "00000001000010000101100000000110";
                        f_reg(114) <= "00000010110101101100100000000110";
                        f_reg(115) <= "00010100110101000000000100110100";
                        f_reg(116) <= "10101100000001100000010010011000";
                        f_reg(117) <= "00000000110010010110000000100000";
                        f_reg(118) <= "00000010100101111101000000100000";
                        f_reg(119) <= "00000001001010000110100000100000";
                        f_reg(120) <= "00000010111101101101100000100000";
                        f_reg(121) <= "00000000001011000111000000000110";
                        f_reg(122) <= "00000001111110101110000000000110";
                        f_reg(123) <= "00000001110010100001000000000110";
                        f_reg(124) <= "00000011100110001000000000000110";
                        f_reg(125) <= "00101001011000110010110110100111";
                        f_reg(126) <= "00101011001100010010110110100111";
                        f_reg(127) <= "00010100001011110000000100101000";
                        f_reg(128) <= "10101100000000010000010010011100";
                        f_reg(129) <= "00000001001001000100000000000110";
                        f_reg(130) <= "00000010111100101011000000000110";
                        f_reg(131) <= "00000000001001110111000000000100";
                        f_reg(132) <= "00000001111101011110000000000100";
                        f_reg(133) <= "00010100110101000000000100100010";
                        f_reg(134) <= "10101100000001100000010010100000";
                        f_reg(135) <= "00000000000000000000000000000000";
                        f_reg(136) <= "00000000000000000000000000000000";
                        f_reg(137) <= "00000000000011000011100101000010";
                        f_reg(138) <= "00000000000110101010100101000010";
                        f_reg(139) <= "00010101100110100000000100011100";
                        f_reg(140) <= "10101100000011000000010011011000";
                        f_reg(141) <= "00000001110001100110000000100010";
                        f_reg(142) <= "00000011100101001101000000100010";
                        f_reg(143) <= "00000001011000110011000000100111";
                        f_reg(144) <= "00000011001100011010000000100111";
                        f_reg(145) <= "00010101101110110000000100010110";
                        f_reg(146) <= "10101100000011010000010010100100";
                        f_reg(147) <= "00000000011010010110100000100100";
                        f_reg(148) <= "00000010001101111101100000100100";
                        f_reg(149) <= "00000000100011100001100000100101";
                        f_reg(150) <= "00000010010111001000100000100101";
                        f_reg(151) <= "00000001000001110100100000100110";
                        f_reg(152) <= "00000010110101011011100000100110";
                        f_reg(153) <= "00111100000001000000101100011101";
                        f_reg(154) <= "00111100000100100000101100011101";
                        f_reg(155) <= "00000000100001110111000000100010";
                        f_reg(156) <= "00000010010101011110000000100010";
                        f_reg(157) <= "00000000000010000011100010000010";
                        f_reg(158) <= "00000000000101101010100010000010";
                        f_reg(159) <= "00000001110011100100000000000100";
                        f_reg(160) <= "00000011100111001011000000000100";
                        f_reg(161) <= "00010100110101000000000100000110";
                        f_reg(162) <= "10101100000001100000010011011100";
                        f_reg(163) <= "00000000000010000011000000100111";
                        f_reg(164) <= "00000000000101101010000000100111";
                        f_reg(165) <= "00010100110101000000000100000010";
                        f_reg(166) <= "10101100000001100000010011100000";
                        f_reg(167) <= "00101101001001101000101000001000";
                        f_reg(168) <= "00101110111101001000101000001000";
                        f_reg(169) <= "00000001101011000100100000100111";
                        f_reg(170) <= "00000011011110101011100000100111";
                        f_reg(171) <= "00010101100110100000000011111100";
                        f_reg(172) <= "10101100000011000000010011100100";
                        f_reg(173) <= "00000000111000100110000000100001";
                        f_reg(174) <= "00000010101100001101000000100001";
                        f_reg(175) <= "00111100000001110011100101100011";
                        f_reg(176) <= "00111100000101010011100101100011";
                        f_reg(177) <= "00000000110001000001000000100111";
                        f_reg(178) <= "00000010100100101000000000100111";
                        f_reg(179) <= "00010100010100000000000011110100";
                        f_reg(180) <= "10101100000000100000010011101000";
                        f_reg(181) <= "00000000000010100001001110000010";
                        f_reg(182) <= "00000000000110001000001110000010";
                        f_reg(183) <= "00000001101000000101000000100000";
                        f_reg(184) <= "00000011011000001100000000100000";
                        f_reg(185) <= "00000000000000000000000000000000";
                        f_reg(186) <= "00000000000000000000000000000000";
                        f_reg(187) <= "00100100100011011111100000101100";
                        f_reg(188) <= "00100110010110111111100000101100";
                        f_reg(189) <= "00101000110001000001110110011111";
                        f_reg(190) <= "00101010100100100001110110011111";
                        f_reg(191) <= "10001100000001100000010011011100";
                        f_reg(192) <= "10001100000101000000010011011100";
                        f_reg(193) <= "00010100110101001111111111111110";
                        f_reg(194) <= "00010101000101100000000011100101";
                        f_reg(195) <= "10101100000010000000010011011100";
                        f_reg(196) <= "00000001110001100100000000100000";
                        f_reg(197) <= "00000011100101001011000000100000";
                        f_reg(198) <= "00000001011000110111000000100001";
                        f_reg(199) <= "00000011001100011110000000100001";
                        f_reg(200) <= "00000001101010000101100000100101";
                        f_reg(201) <= "00000011011101101100100000100101";
                        f_reg(202) <= "00000000010001110001100000000111";
                        f_reg(203) <= "00000010000101011000100000000111";
                        f_reg(204) <= "00000001001011000110100000100001";
                        f_reg(205) <= "00000010111110101101100000100001";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101100001000010001100101111000";
                        f_reg(209) <= "00101101111011110001100101111000";
                        f_reg(210) <= "00010101010110000000000011010101";
                        f_reg(211) <= "10101100000010100000010010101000";
                        f_reg(212) <= "00000001011001010100000000100100";
                        f_reg(213) <= "00000011001100111011000000100100";
                        f_reg(214) <= "00010101000101100000000011010001";
                        f_reg(215) <= "10101100000010000000010010101100";
                        f_reg(216) <= "10001100000001110000010011011100";
                        f_reg(217) <= "10001100000101010000010011011100";
                        f_reg(218) <= "00010100111101011111111111111110";
                        f_reg(219) <= "00000000111001000001000000100000";
                        f_reg(220) <= "00000010101100101000000000100000";
                        f_reg(221) <= "00000000010001100100100000100000";
                        f_reg(222) <= "00000010000101001011100000100000";
                        f_reg(223) <= "00000000000001100110011011000011";
                        f_reg(224) <= "00000000000101001101011011000011";
                        f_reg(225) <= "00000001110011000110000000000100";
                        f_reg(226) <= "00000011100110101101000000000100";
                        f_reg(227) <= "10001100000010100000010011100100";
                        f_reg(228) <= "10001100000110000000010011100100";
                        f_reg(229) <= "00010101010110001111111111111110";
                        f_reg(230) <= "10001100000010110000010011011000";
                        f_reg(231) <= "10001100000110010000010011011000";
                        f_reg(232) <= "00010101011110011111111111111110";
                        f_reg(233) <= "00000001010010110010100000101010";
                        f_reg(234) <= "00000011000110011001100000101010";
                        f_reg(235) <= "10001100000010000000010011100000";
                        f_reg(236) <= "10001100000101100000010011100000";
                        f_reg(237) <= "00010101000101101111111111111110";
                        f_reg(238) <= "00000001000011010011100000101011";
                        f_reg(239) <= "00000010110110111010100000101011";
                        f_reg(240) <= "00010100110101000000000010110111";
                        f_reg(241) <= "10101100000001100000010010110000";
                        f_reg(242) <= "00110001100001001010010100111111";
                        f_reg(243) <= "00110011010100101010010100111111";
                        f_reg(244) <= "10001100000000100000010011101000";
                        f_reg(245) <= "10001100000100000000010011101000";
                        f_reg(246) <= "00010100010100001111111111111110";
                        f_reg(247) <= "00000000011000100111000000000110";
                        f_reg(248) <= "00000010001100001110000000000110";
                        f_reg(249) <= "00000000111001010101000000100111";
                        f_reg(250) <= "00000010101100111100000000100111";
                        f_reg(251) <= "00100001010010111101011101010111";
                        f_reg(252) <= "00100011000110011101011101010111";
                        f_reg(253) <= "00101000100010000001110011001011";
                        f_reg(254) <= "00101010010101100001110011001011";
                        f_reg(255) <= "00010101110111000000000010101000";
                        f_reg(256) <= "10101100000011100000010010110100";
                        f_reg(257) <= "00010100101100110000000010100110";
                        f_reg(258) <= "10101100000001010000010010111000";
                        f_reg(259) <= "00010101001101110000000010100100";
                        f_reg(260) <= "10101100000010010000010010111100";
                        f_reg(261) <= "00010101110111000000000010100010";
                        f_reg(262) <= "10101100000011100000010011000000";
                        f_reg(263) <= "00111000111011011011111110101011";
                        f_reg(264) <= "00111010101110111011111110101011";
                        f_reg(265) <= "00101001011001101011000111001110";
                        f_reg(266) <= "00101011001101001011000111001110";
                        f_reg(267) <= "00010100001011110000000010011100";
                        f_reg(268) <= "10101100000000010000010011000100";
                        f_reg(269) <= "00010100110101000000000010011010";
                        f_reg(270) <= "10101100000001100000010011001000";
                        f_reg(271) <= "00100001101011000011010101111100";
                        f_reg(272) <= "00100011011110100011010101111100";
                        f_reg(273) <= "00010100011100010000000010010110";
                        f_reg(274) <= "10101100000000110000010011001100";
                        f_reg(275) <= "00000001100010110001000000100100";
                        f_reg(276) <= "00000011010110011000000000100100";
                        f_reg(277) <= "00100000010010100001001001100010";
                        f_reg(278) <= "00100010000110000001001001100010";
                        f_reg(279) <= "00010101000101100000000010010000";
                        f_reg(280) <= "10101100000010000000010011010000";
                        f_reg(281) <= "00010101010110000000000010001110";
                        f_reg(282) <= "10101100000010100000010011010100";
                        f_reg(283) <= "00100011110111011111111100000110";
                        f_reg(284) <= "00010011101000000000000000100000";
                        f_reg(285) <= "00100011110111011111111000001100";
                        f_reg(286) <= "00010011101000000000000000011110";
                        f_reg(287) <= "00100011110111011111110100010010";
                        f_reg(288) <= "00010011101000000000000000011100";
                        f_reg(289) <= "00100011110111101111111111111111";
                        f_reg(290) <= "00100011111111111111111111111111";
                        f_reg(291) <= "00010111110111110000000010000100";
                        f_reg(292) <= "00011111111000001111111100110111";
                        f_reg(293) <= "00010000000000000000000100001111";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "00000000000000000000000000000000";
                        f_reg(304) <= "00000000000000000000000000000000";
                        f_reg(305) <= "00000000000000000000000000000000";
                        f_reg(306) <= "00000000000000000000000000000000";
                        f_reg(307) <= "00000000000000000000000000000000";
                        f_reg(308) <= "00000000000000000000000000000000";
                        f_reg(309) <= "00000000000000000000000000000000";
                        f_reg(310) <= "00000000000000000000000000000000";
                        f_reg(311) <= "00000000000000000000000000000000";
                        f_reg(312) <= "00000000000000000000000000000000";
                        f_reg(313) <= "00000000000000000000000000000000";
                        f_reg(314) <= "00000000000000000000000000000000";
                        f_reg(315) <= "00000000000000000000000000000000";
                        f_reg(316) <= "10001100000111010000100001000000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010100001011110000000001100110";
                        f_reg(322) <= "10101111101000010000011111001000";
                        f_reg(323) <= "10001100000111010000100001000000";
                        f_reg(324) <= "00011111101000000000000000000011";
                        f_reg(325) <= "00100000000111010000000000111100";
                        f_reg(326) <= "00010000000000000000000000000010";
                        f_reg(327) <= "00100000000111010000000000000000";
                        f_reg(328) <= "00010100010100000000000001011111";
                        f_reg(329) <= "10101111101000100000011111001100";
                        f_reg(330) <= "10001100000111010000100001000000";
                        f_reg(331) <= "00011111101000000000000000000011";
                        f_reg(332) <= "00100000000111010000000000111100";
                        f_reg(333) <= "00010000000000000000000000000010";
                        f_reg(334) <= "00100000000111010000000000000000";
                        f_reg(335) <= "00010100011100010000000001011000";
                        f_reg(336) <= "10101111101000110000011111010000";
                        f_reg(337) <= "10001100000111010000100001000000";
                        f_reg(338) <= "00011111101000000000000000000011";
                        f_reg(339) <= "00100000000111010000000000111100";
                        f_reg(340) <= "00010000000000000000000000000010";
                        f_reg(341) <= "00100000000111010000000000000000";
                        f_reg(342) <= "00010100100100100000000001010001";
                        f_reg(343) <= "10101111101001000000011111010100";
                        f_reg(344) <= "10001100000111010000100001000000";
                        f_reg(345) <= "00011111101000000000000000000011";
                        f_reg(346) <= "00100000000111010000000000111100";
                        f_reg(347) <= "00010000000000000000000000000010";
                        f_reg(348) <= "00100000000111010000000000000000";
                        f_reg(349) <= "00010100101100110000000001001010";
                        f_reg(350) <= "10101111101001010000011111011000";
                        f_reg(351) <= "10001100000111010000100001000000";
                        f_reg(352) <= "00011111101000000000000000000011";
                        f_reg(353) <= "00100000000111010000000000111100";
                        f_reg(354) <= "00010000000000000000000000000010";
                        f_reg(355) <= "00100000000111010000000000000000";
                        f_reg(356) <= "00010100110101000000000001000011";
                        f_reg(357) <= "10101111101001100000011111011100";
                        f_reg(358) <= "10001100000111010000100001000000";
                        f_reg(359) <= "00011111101000000000000000000011";
                        f_reg(360) <= "00100000000111010000000000111100";
                        f_reg(361) <= "00010000000000000000000000000010";
                        f_reg(362) <= "00100000000111010000000000000000";
                        f_reg(363) <= "00010100111101010000000000111100";
                        f_reg(364) <= "10101111101001110000011111100000";
                        f_reg(365) <= "10001100000111010000100001000000";
                        f_reg(366) <= "00011111101000000000000000000011";
                        f_reg(367) <= "00100000000111010000000000111100";
                        f_reg(368) <= "00010000000000000000000000000010";
                        f_reg(369) <= "00100000000111010000000000000000";
                        f_reg(370) <= "00010101000101100000000000110101";
                        f_reg(371) <= "10101111101010000000011111100100";
                        f_reg(372) <= "10001100000111010000100001000000";
                        f_reg(373) <= "00011111101000000000000000000011";
                        f_reg(374) <= "00100000000111010000000000111100";
                        f_reg(375) <= "00010000000000000000000000000010";
                        f_reg(376) <= "00100000000111010000000000000000";
                        f_reg(377) <= "00010101001101110000000000101110";
                        f_reg(378) <= "10101111101010010000011111101000";
                        f_reg(379) <= "10001100000111010000100001000000";
                        f_reg(380) <= "00011111101000000000000000000011";
                        f_reg(381) <= "00100000000111010000000000111100";
                        f_reg(382) <= "00010000000000000000000000000010";
                        f_reg(383) <= "00100000000111010000000000000000";
                        f_reg(384) <= "00010101010110000000000000100111";
                        f_reg(385) <= "10101111101010100000011111101100";
                        f_reg(386) <= "10001100000111010000100001000000";
                        f_reg(387) <= "00011111101000000000000000000011";
                        f_reg(388) <= "00100000000111010000000000111100";
                        f_reg(389) <= "00010000000000000000000000000010";
                        f_reg(390) <= "00100000000111010000000000000000";
                        f_reg(391) <= "00010101011110010000000000100000";
                        f_reg(392) <= "10101111101010110000011111110000";
                        f_reg(393) <= "10001100000111010000100001000000";
                        f_reg(394) <= "00011111101000000000000000000011";
                        f_reg(395) <= "00100000000111010000000000111100";
                        f_reg(396) <= "00010000000000000000000000000010";
                        f_reg(397) <= "00100000000111010000000000000000";
                        f_reg(398) <= "00010101100110100000000000011001";
                        f_reg(399) <= "10101111101011000000011111110100";
                        f_reg(400) <= "10001100000111010000100001000000";
                        f_reg(401) <= "00011111101000000000000000000011";
                        f_reg(402) <= "00100000000111010000000000111100";
                        f_reg(403) <= "00010000000000000000000000000010";
                        f_reg(404) <= "00100000000111010000000000000000";
                        f_reg(405) <= "00010101101110110000000000010010";
                        f_reg(406) <= "10101111101011010000011111111000";
                        f_reg(407) <= "10001100000111010000100001000000";
                        f_reg(408) <= "00011111101000000000000000000011";
                        f_reg(409) <= "00100000000111010000000000111100";
                        f_reg(410) <= "00010000000000000000000000000010";
                        f_reg(411) <= "00100000000111010000000000000000";
                        f_reg(412) <= "00010101110111000000000000001011";
                        f_reg(413) <= "10101111101011100000011111111100";
                        f_reg(414) <= "10001100000111010000100001000000";
                        f_reg(415) <= "00011111101000000000000000000011";
                        f_reg(416) <= "00100000000111010000000000111100";
                        f_reg(417) <= "00010000000000000000000000000010";
                        f_reg(418) <= "00100000000111010000000000000000";
                        f_reg(419) <= "00010111110111110000000000000100";
                        f_reg(420) <= "10101111101111100000100000000000";
                        f_reg(421) <= "10101100000111010000100001000000";
                        f_reg(422) <= "00010000000000001111111101111011";
                        f_reg(423) <= "10001100000111010000100001000000";
                        f_reg(424) <= "10001111101000010000011111001000";
                        f_reg(425) <= "10001100000111010000100001000000";
                        f_reg(426) <= "10001111101011110000011111001000";
                        f_reg(427) <= "00010100001011111111111111111100";
                        f_reg(428) <= "10001100000111010000100001000000";
                        f_reg(429) <= "10001111101000100000011111001100";
                        f_reg(430) <= "10001100000111010000100001000000";
                        f_reg(431) <= "10001111101100000000011111001100";
                        f_reg(432) <= "00010100010100001111111111111100";
                        f_reg(433) <= "10001100000111010000100001000000";
                        f_reg(434) <= "10001111101000110000011111010000";
                        f_reg(435) <= "10001100000111010000100001000000";
                        f_reg(436) <= "10001111101100010000011111010000";
                        f_reg(437) <= "00010100011100011111111111111100";
                        f_reg(438) <= "10001100000111010000100001000000";
                        f_reg(439) <= "10001111101001000000011111010100";
                        f_reg(440) <= "10001100000111010000100001000000";
                        f_reg(441) <= "10001111101100100000011111010100";
                        f_reg(442) <= "00010100100100101111111111111100";
                        f_reg(443) <= "10001100000111010000100001000000";
                        f_reg(444) <= "10001111101001010000011111011000";
                        f_reg(445) <= "10001100000111010000100001000000";
                        f_reg(446) <= "10001111101100110000011111011000";
                        f_reg(447) <= "00010100101100111111111111111100";
                        f_reg(448) <= "10001100000111010000100001000000";
                        f_reg(449) <= "10001111101001100000011111011100";
                        f_reg(450) <= "10001100000111010000100001000000";
                        f_reg(451) <= "10001111101101000000011111011100";
                        f_reg(452) <= "00010100110101001111111111111100";
                        f_reg(453) <= "10001100000111010000100001000000";
                        f_reg(454) <= "10001111101001110000011111100000";
                        f_reg(455) <= "10001100000111010000100001000000";
                        f_reg(456) <= "10001111101101010000011111100000";
                        f_reg(457) <= "00010100111101011111111111111100";
                        f_reg(458) <= "10001100000111010000100001000000";
                        f_reg(459) <= "10001111101010000000011111100100";
                        f_reg(460) <= "10001100000111010000100001000000";
                        f_reg(461) <= "10001111101101100000011111100100";
                        f_reg(462) <= "00010101000101101111111111111100";
                        f_reg(463) <= "10001100000111010000100001000000";
                        f_reg(464) <= "10001111101010010000011111101000";
                        f_reg(465) <= "10001100000111010000100001000000";
                        f_reg(466) <= "10001111101101110000011111101000";
                        f_reg(467) <= "00010101001101111111111111111100";
                        f_reg(468) <= "10001100000111010000100001000000";
                        f_reg(469) <= "10001111101010100000011111101100";
                        f_reg(470) <= "10001100000111010000100001000000";
                        f_reg(471) <= "10001111101110000000011111101100";
                        f_reg(472) <= "00010101010110001111111111111100";
                        f_reg(473) <= "10001100000111010000100001000000";
                        f_reg(474) <= "10001111101010110000011111110000";
                        f_reg(475) <= "10001100000111010000100001000000";
                        f_reg(476) <= "10001111101110010000011111110000";
                        f_reg(477) <= "00010101011110011111111111111100";
                        f_reg(478) <= "10001100000111010000100001000000";
                        f_reg(479) <= "10001111101011000000011111110100";
                        f_reg(480) <= "10001100000111010000100001000000";
                        f_reg(481) <= "10001111101110100000011111110100";
                        f_reg(482) <= "00010101100110101111111111111100";
                        f_reg(483) <= "10001100000111010000100001000000";
                        f_reg(484) <= "10001111101011010000011111111000";
                        f_reg(485) <= "10001100000111010000100001000000";
                        f_reg(486) <= "10001111101110110000011111111000";
                        f_reg(487) <= "00010101101110111111111111111100";
                        f_reg(488) <= "10001100000111010000100001000000";
                        f_reg(489) <= "10001111101011100000011111111100";
                        f_reg(490) <= "10001100000111010000100001000000";
                        f_reg(491) <= "10001111101111000000011111111100";
                        f_reg(492) <= "00010101110111001111111111111100";
                        f_reg(493) <= "10001100000111010000100001000000";
                        f_reg(494) <= "10001111101111100000100000000000";
                        f_reg(495) <= "10001100000111010000100001000000";
                        f_reg(496) <= "10001111101111110000100000000000";
                        f_reg(497) <= "00010111110111111111111111111100";
                        f_reg(498) <= "00010000000000001111111100101111";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000001111100111";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                        f_reg(551) <= "00000000000000000000000000000000";
                        f_reg(552) <= "00000000000000000000000000000000";
                        f_reg(553) <= "00000000000000000000000000000000";
                        f_reg(554) <= "00000000000000000000000000000000";
                        f_reg(555) <= "00000000000000000000000000000000";
                        f_reg(556) <= "00000000000000000000000000000000";
                        f_reg(557) <= "00000000000000000000000000000000";
                        f_reg(558) <= "00000000000000000000000000000000";
                        f_reg(559) <= "00000000000000000000000000000000";
                        f_reg(560) <= "00000000000000000000000000000000";
                        f_reg(561) <= "00000000000000000000000000000000";
                        f_reg(562) <= "00000000000000000000000000000000";
                        f_reg(563) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010000111101001010";
                        f_reg(4) <= "00111000000000101100101100111110";
                        f_reg(5) <= "10101100000000010000010010010100";
                        f_reg(6) <= "00000000000000000001110100000010";
                        f_reg(7) <= "00000000001000100010000000100011";
                        f_reg(8) <= "00111000010001010010110011000011";
                        f_reg(9) <= "00110000100001100101101111111001";
                        f_reg(10) <= "00000000010001100011100000100000";
                        f_reg(11) <= "00000000011000100100000000100010";
                        f_reg(12) <= "00100100100010011101110001100011";
                        f_reg(13) <= "00110000011010100001111000100100";
                        f_reg(14) <= "00000001000010000101100000000110";
                        f_reg(15) <= "10101100000001100000010010011000";
                        f_reg(16) <= "00000000110010010110000000100000";
                        f_reg(17) <= "00000001001010000110100000100000";
                        f_reg(18) <= "00000000001011000111000000000110";
                        f_reg(19) <= "00000001110010100111100000000110";
                        f_reg(20) <= "00101001011100000010110110100111";
                        f_reg(21) <= "10101100000000010000010010011100";
                        f_reg(22) <= "00000001001001001000100000000110";
                        f_reg(23) <= "00000000001001111001000000000100";
                        f_reg(24) <= "10101100000001100000010010100000";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00000000000011001001100101000010";
                        f_reg(27) <= "00000010010001101010000000100010";
                        f_reg(28) <= "00000001011100001010100000100111";
                        f_reg(29) <= "10101100000011010000010010100100";
                        f_reg(30) <= "00000010000010011011000000100100";
                        f_reg(31) <= "00000000100100101011100000100101";
                        f_reg(32) <= "00000010001100111100000000100110";
                        f_reg(33) <= "00111100000110010000101100011101";
                        f_reg(34) <= "00000011001100111101000000100010";
                        f_reg(35) <= "00000000000100011101100010000010";
                        f_reg(36) <= "00000011010110101110000000000100";
                        f_reg(37) <= "00000000000111001110100000100111";
                        f_reg(38) <= "00101111000111101000101000001000";
                        f_reg(39) <= "00000010110101000001000000100111";
                        f_reg(40) <= "00000011011011110001100000100001";
                        f_reg(41) <= "00111100000010000011100101100011";
                        f_reg(42) <= "00000011110110010111000000100111";
                        f_reg(43) <= "00000000000010100011101110000010";
                        f_reg(44) <= "00000010110000000011000000100000";
                        f_reg(45) <= "00000000000000000000000000000000";
                        f_reg(46) <= "00100111001011011111100000101100";
                        f_reg(47) <= "00101011110100000001110110011111";
                        f_reg(48) <= "00000011010101010100100000100000";
                        f_reg(49) <= "00000001011101110010000000100001";
                        f_reg(50) <= "00000001101010011001000000100101";
                        f_reg(51) <= "00000000111010001001100000000111";
                        f_reg(52) <= "00000000010000111000100000100001";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00101100001000010001100101111000";
                        f_reg(55) <= "10101100000001100000010010101000";
                        f_reg(56) <= "00000010010001011100000000100100";
                        f_reg(57) <= "10101100000110000000010010101100";
                        f_reg(58) <= "00000011100100001101100000100000";
                        f_reg(59) <= "00000011011101010111100000100000";
                        f_reg(60) <= "00000000000101010101011011000011";
                        f_reg(61) <= "00000000100010100101000000000100";
                        f_reg(62) <= "00000010100011001011000000101010";
                        f_reg(63) <= "00000011101100011100100000101011";
                        f_reg(64) <= "10101100000101010000010010110000";
                        f_reg(65) <= "00110001010111101010010100111111";
                        f_reg(66) <= "00000010011011101101000000000110";
                        f_reg(67) <= "00000011001101100101100000100111";
                        f_reg(68) <= "00100001011101111101011101010111";
                        f_reg(69) <= "00101011110011010001110011001011";
                        f_reg(70) <= "10101100000110100000010010110100";
                        f_reg(71) <= "10101100000101100000010010111000";
                        f_reg(72) <= "10101100000011110000010010111100";
                        f_reg(73) <= "10101100000110100000010011000000";
                        f_reg(74) <= "00111011001010011011111110101011";
                        f_reg(75) <= "00101010111010001011000111001110";
                        f_reg(76) <= "10101100000000010000010011000100";
                        f_reg(77) <= "10101100000010000000010011001000";
                        f_reg(78) <= "00100001001001110011010101111100";
                        f_reg(79) <= "10101100000100110000010011001100";
                        f_reg(80) <= "00000000111101110001000000100100";
                        f_reg(81) <= "00100000010000110001001001100010";
                        f_reg(82) <= "10101100000011010000010011010000";
                        f_reg(83) <= "10101100000000110000010011010100";
                        f_reg(84) <= "00100011111111111111111111111111";
                        f_reg(85) <= "00011111111000001111111110101110";
                        f_reg(86) <= "00010000000000000000000111011110";
                        f_reg(87) <= "00111100000111100000001111100111";
                        f_reg(88) <= "00111100000111110000001111100111";
                        f_reg(89) <= "00000000000111101111010000000010";
                        f_reg(90) <= "00000000000111111111110000000010";
                        f_reg(91) <= "00111100000000010000111101001010";
                        f_reg(92) <= "00111100000011110000111101001010";
                        f_reg(93) <= "00111000000000101100101100111110";
                        f_reg(94) <= "00111000000100001100101100111110";
                        f_reg(95) <= "00010100001011110000000101001000";
                        f_reg(96) <= "10101100000000010000010010010100";
                        f_reg(97) <= "00000000000000000001110100000010";
                        f_reg(98) <= "00000000000000001000110100000010";
                        f_reg(99) <= "00000000001000100010000000100011";
                        f_reg(100) <= "00000001111100001001000000100011";
                        f_reg(101) <= "00111000010001010010110011000011";
                        f_reg(102) <= "00111010000100110010110011000011";
                        f_reg(103) <= "00110000100001100101101111111001";
                        f_reg(104) <= "00110010010101000101101111111001";
                        f_reg(105) <= "00000000010001100011100000100000";
                        f_reg(106) <= "00000010000101001010100000100000";
                        f_reg(107) <= "00000000011000100100000000100010";
                        f_reg(108) <= "00000010001100001011000000100010";
                        f_reg(109) <= "00100100100010011101110001100011";
                        f_reg(110) <= "00100110010101111101110001100011";
                        f_reg(111) <= "00110000011010100001111000100100";
                        f_reg(112) <= "00110010001110000001111000100100";
                        f_reg(113) <= "00000001000010000101100000000110";
                        f_reg(114) <= "00000010110101101100100000000110";
                        f_reg(115) <= "00010100110101000000000100110100";
                        f_reg(116) <= "10101100000001100000010010011000";
                        f_reg(117) <= "00000000110010010110000000100000";
                        f_reg(118) <= "00000010100101111101000000100000";
                        f_reg(119) <= "00000001001010000110100000100000";
                        f_reg(120) <= "00000010111101101101100000100000";
                        f_reg(121) <= "00000000001011000111000000000110";
                        f_reg(122) <= "00000001111110101110000000000110";
                        f_reg(123) <= "00000001110010100001000000000110";
                        f_reg(124) <= "00000011100110001000000000000110";
                        f_reg(125) <= "00101001011000110010110110100111";
                        f_reg(126) <= "00101011001100010010110110100111";
                        f_reg(127) <= "00010100001011110000000100101000";
                        f_reg(128) <= "10101100000000010000010010011100";
                        f_reg(129) <= "00000001001001000100000000000110";
                        f_reg(130) <= "00000010111100101011000000000110";
                        f_reg(131) <= "00000000001001110111000000000100";
                        f_reg(132) <= "00000001111101011110000000000100";
                        f_reg(133) <= "00010100110101000000000100100010";
                        f_reg(134) <= "10101100000001100000010010100000";
                        f_reg(135) <= "00000000000000000000000000000000";
                        f_reg(136) <= "00000000000000000000000000000000";
                        f_reg(137) <= "00000000000011000011100101000010";
                        f_reg(138) <= "00000000000110101010100101000010";
                        f_reg(139) <= "00010101100110100000000100011100";
                        f_reg(140) <= "10101100000011000000010011011000";
                        f_reg(141) <= "00000001110001100110000000100010";
                        f_reg(142) <= "00000011100101001101000000100010";
                        f_reg(143) <= "00000001011000110011000000100111";
                        f_reg(144) <= "00000011001100011010000000100111";
                        f_reg(145) <= "00010101101110110000000100010110";
                        f_reg(146) <= "10101100000011010000010010100100";
                        f_reg(147) <= "00000000011010010110100000100100";
                        f_reg(148) <= "00000010001101111101100000100100";
                        f_reg(149) <= "00000000100011100001100000100101";
                        f_reg(150) <= "00000010010111001000100000100101";
                        f_reg(151) <= "00000001000001110100100000100110";
                        f_reg(152) <= "00000010110101011011100000100110";
                        f_reg(153) <= "00111100000001000000101100011101";
                        f_reg(154) <= "00111100000100100000101100011101";
                        f_reg(155) <= "00000000100001110111000000100010";
                        f_reg(156) <= "00000010010101011110000000100010";
                        f_reg(157) <= "00000000000010000011100010000010";
                        f_reg(158) <= "00000000000101101010100010000010";
                        f_reg(159) <= "00000001110011100100000000000100";
                        f_reg(160) <= "00000011100111001011000000000100";
                        f_reg(161) <= "00010100110101000000000100000110";
                        f_reg(162) <= "10101100000001100000010011011100";
                        f_reg(163) <= "00000000000010000011000000100111";
                        f_reg(164) <= "00000000000101101010000000100111";
                        f_reg(165) <= "00010100110101000000000100000010";
                        f_reg(166) <= "10101100000001100000010011100000";
                        f_reg(167) <= "00101101001001101000101000001000";
                        f_reg(168) <= "00101110111101001000101000001000";
                        f_reg(169) <= "00000001101011000100100000100111";
                        f_reg(170) <= "00000011011110101011100000100111";
                        f_reg(171) <= "00010101100110100000000011111100";
                        f_reg(172) <= "10101100000011000000010011100100";
                        f_reg(173) <= "00000000111000100110000000100001";
                        f_reg(174) <= "00000010101100001101000000100001";
                        f_reg(175) <= "00111100000001110011100101100011";
                        f_reg(176) <= "00111100000101010011100101100011";
                        f_reg(177) <= "00000000110001000001000000100111";
                        f_reg(178) <= "00000010100100101000000000100111";
                        f_reg(179) <= "00010100010100000000000011110100";
                        f_reg(180) <= "10101100000000100000010011101000";
                        f_reg(181) <= "00000000000010100001001110000010";
                        f_reg(182) <= "00000000000110001000001110000010";
                        f_reg(183) <= "00000001101000000101000000100000";
                        f_reg(184) <= "00000011011000001100000000100000";
                        f_reg(185) <= "00000000000000000000000000000000";
                        f_reg(186) <= "00000000000000000000000000000000";
                        f_reg(187) <= "00100100100011011111100000101100";
                        f_reg(188) <= "00100110010110111111100000101100";
                        f_reg(189) <= "00101000110001000001110110011111";
                        f_reg(190) <= "00101010100100100001110110011111";
                        f_reg(191) <= "10001100000001100000010011011100";
                        f_reg(192) <= "10001100000101000000010011011100";
                        f_reg(193) <= "00010100110101001111111111111110";
                        f_reg(194) <= "00010101000101100000000011100101";
                        f_reg(195) <= "10101100000010000000010011011100";
                        f_reg(196) <= "00000001110001100100000000100000";
                        f_reg(197) <= "00000011100101001011000000100000";
                        f_reg(198) <= "00000001011000110111000000100001";
                        f_reg(199) <= "00000011001100011110000000100001";
                        f_reg(200) <= "00000001101010000101100000100101";
                        f_reg(201) <= "00000011011101101100100000100101";
                        f_reg(202) <= "00000000010001110001100000000111";
                        f_reg(203) <= "00000010000101011000100000000111";
                        f_reg(204) <= "00000001001011000110100000100001";
                        f_reg(205) <= "00000010111110101101100000100001";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101100001000010001100101111000";
                        f_reg(209) <= "00101101111011110001100101111000";
                        f_reg(210) <= "00010101010110000000000011010101";
                        f_reg(211) <= "10101100000010100000010010101000";
                        f_reg(212) <= "00000001011001010100000000100100";
                        f_reg(213) <= "00000011001100111011000000100100";
                        f_reg(214) <= "00010101000101100000000011010001";
                        f_reg(215) <= "10101100000010000000010010101100";
                        f_reg(216) <= "10001100000001110000010011011100";
                        f_reg(217) <= "10001100000101010000010011011100";
                        f_reg(218) <= "00010100111101011111111111111110";
                        f_reg(219) <= "00000000111001000001000000100000";
                        f_reg(220) <= "00000010101100101000000000100000";
                        f_reg(221) <= "00000000010001100100100000100000";
                        f_reg(222) <= "00000010000101001011100000100000";
                        f_reg(223) <= "00000000000001100110011011000011";
                        f_reg(224) <= "00000000000101001101011011000011";
                        f_reg(225) <= "00000001110011000110000000000100";
                        f_reg(226) <= "00000011100110101101000000000100";
                        f_reg(227) <= "10001100000010100000010011100100";
                        f_reg(228) <= "10001100000110000000010011100100";
                        f_reg(229) <= "00010101010110001111111111111110";
                        f_reg(230) <= "10001100000010110000010011011000";
                        f_reg(231) <= "10001100000110010000010011011000";
                        f_reg(232) <= "00010101011110011111111111111110";
                        f_reg(233) <= "00000001010010110010100000101010";
                        f_reg(234) <= "00000011000110011001100000101010";
                        f_reg(235) <= "10001100000010000000010011100000";
                        f_reg(236) <= "10001100000101100000010011100000";
                        f_reg(237) <= "00010101000101101111111111111110";
                        f_reg(238) <= "00000001000011010011100000101011";
                        f_reg(239) <= "00000010110110111010100000101011";
                        f_reg(240) <= "00010100110101000000000010110111";
                        f_reg(241) <= "10101100000001100000010010110000";
                        f_reg(242) <= "00110001100001001010010100111111";
                        f_reg(243) <= "00110011010100101010010100111111";
                        f_reg(244) <= "10001100000000100000010011101000";
                        f_reg(245) <= "10001100000100000000010011101000";
                        f_reg(246) <= "00010100010100001111111111111110";
                        f_reg(247) <= "00000000011000100111000000000110";
                        f_reg(248) <= "00000010001100001110000000000110";
                        f_reg(249) <= "00000000111001010101000000100111";
                        f_reg(250) <= "00000010101100111100000000100111";
                        f_reg(251) <= "00100001010010111101011101010111";
                        f_reg(252) <= "00100011000110011101011101010111";
                        f_reg(253) <= "00101000100010000001110011001011";
                        f_reg(254) <= "00101010010101100001110011001011";
                        f_reg(255) <= "00010101110111000000000010101000";
                        f_reg(256) <= "10101100000011100000010010110100";
                        f_reg(257) <= "00010100101100110000000010100110";
                        f_reg(258) <= "10101100000001010000010010111000";
                        f_reg(259) <= "00010101001101110000000010100100";
                        f_reg(260) <= "10101100000010010000010010111100";
                        f_reg(261) <= "00010101110111000000000010100010";
                        f_reg(262) <= "10101100000011100000010011000000";
                        f_reg(263) <= "00111000111011011011111110101011";
                        f_reg(264) <= "00111010101110111011111110101011";
                        f_reg(265) <= "00101001011001101011000111001110";
                        f_reg(266) <= "00101011001101001011000111001110";
                        f_reg(267) <= "00010100001011110000000010011100";
                        f_reg(268) <= "10101100000000010000010011000100";
                        f_reg(269) <= "00010100110101000000000010011010";
                        f_reg(270) <= "10101100000001100000010011001000";
                        f_reg(271) <= "00100001101011000011010101111100";
                        f_reg(272) <= "00100011011110100011010101111100";
                        f_reg(273) <= "00010100011100010000000010010110";
                        f_reg(274) <= "10101100000000110000010011001100";
                        f_reg(275) <= "00000001100010110001000000100100";
                        f_reg(276) <= "00000011010110011000000000100100";
                        f_reg(277) <= "00100000010010100001001001100010";
                        f_reg(278) <= "00100010000110000001001001100010";
                        f_reg(279) <= "00010101000101100000000010010000";
                        f_reg(280) <= "10101100000010000000010011010000";
                        f_reg(281) <= "00010101010110000000000010001110";
                        f_reg(282) <= "10101100000010100000010011010100";
                        f_reg(283) <= "00100011110111011111111100000110";
                        f_reg(284) <= "00010011101000000000000000100000";
                        f_reg(285) <= "00100011110111011111111000001100";
                        f_reg(286) <= "00010011101000000000000000011110";
                        f_reg(287) <= "00100011110111011111110100010010";
                        f_reg(288) <= "00010011101000000000000000011100";
                        f_reg(289) <= "00100011110111101111111111111111";
                        f_reg(290) <= "00100011111111111111111111111111";
                        f_reg(291) <= "00010111110111110000000010000100";
                        f_reg(292) <= "00011111111000001111111100110111";
                        f_reg(293) <= "00010000000000000000000100001111";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "00000000000000000000000000000000";
                        f_reg(304) <= "00000000000000000000000000000000";
                        f_reg(305) <= "00000000000000000000000000000000";
                        f_reg(306) <= "00000000000000000000000000000000";
                        f_reg(307) <= "00000000000000000000000000000000";
                        f_reg(308) <= "00000000000000000000000000000000";
                        f_reg(309) <= "00000000000000000000000000000000";
                        f_reg(310) <= "00000000000000000000000000000000";
                        f_reg(311) <= "00000000000000000000000000000000";
                        f_reg(312) <= "00000000000000000000000000000000";
                        f_reg(313) <= "00000000000000000000000000000000";
                        f_reg(314) <= "00000000000000000000000000000000";
                        f_reg(315) <= "00000000000000000000000000000000";
                        f_reg(316) <= "10001100000111010000100001000000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010100001011110000000001100110";
                        f_reg(322) <= "10101111101000010000011111001000";
                        f_reg(323) <= "10001100000111010000100001000000";
                        f_reg(324) <= "00011111101000000000000000000011";
                        f_reg(325) <= "00100000000111010000000000111100";
                        f_reg(326) <= "00010000000000000000000000000010";
                        f_reg(327) <= "00100000000111010000000000000000";
                        f_reg(328) <= "00010100010100000000000001011111";
                        f_reg(329) <= "10101111101000100000011111001100";
                        f_reg(330) <= "10001100000111010000100001000000";
                        f_reg(331) <= "00011111101000000000000000000011";
                        f_reg(332) <= "00100000000111010000000000111100";
                        f_reg(333) <= "00010000000000000000000000000010";
                        f_reg(334) <= "00100000000111010000000000000000";
                        f_reg(335) <= "00010100011100010000000001011000";
                        f_reg(336) <= "10101111101000110000011111010000";
                        f_reg(337) <= "10001100000111010000100001000000";
                        f_reg(338) <= "00011111101000000000000000000011";
                        f_reg(339) <= "00100000000111010000000000111100";
                        f_reg(340) <= "00010000000000000000000000000010";
                        f_reg(341) <= "00100000000111010000000000000000";
                        f_reg(342) <= "00010100100100100000000001010001";
                        f_reg(343) <= "10101111101001000000011111010100";
                        f_reg(344) <= "10001100000111010000100001000000";
                        f_reg(345) <= "00011111101000000000000000000011";
                        f_reg(346) <= "00100000000111010000000000111100";
                        f_reg(347) <= "00010000000000000000000000000010";
                        f_reg(348) <= "00100000000111010000000000000000";
                        f_reg(349) <= "00010100101100110000000001001010";
                        f_reg(350) <= "10101111101001010000011111011000";
                        f_reg(351) <= "10001100000111010000100001000000";
                        f_reg(352) <= "00011111101000000000000000000011";
                        f_reg(353) <= "00100000000111010000000000111100";
                        f_reg(354) <= "00010000000000000000000000000010";
                        f_reg(355) <= "00100000000111010000000000000000";
                        f_reg(356) <= "00010100110101000000000001000011";
                        f_reg(357) <= "10101111101001100000011111011100";
                        f_reg(358) <= "10001100000111010000100001000000";
                        f_reg(359) <= "00011111101000000000000000000011";
                        f_reg(360) <= "00100000000111010000000000111100";
                        f_reg(361) <= "00010000000000000000000000000010";
                        f_reg(362) <= "00100000000111010000000000000000";
                        f_reg(363) <= "00010100111101010000000000111100";
                        f_reg(364) <= "10101111101001110000011111100000";
                        f_reg(365) <= "10001100000111010000100001000000";
                        f_reg(366) <= "00011111101000000000000000000011";
                        f_reg(367) <= "00100000000111010000000000111100";
                        f_reg(368) <= "00010000000000000000000000000010";
                        f_reg(369) <= "00100000000111010000000000000000";
                        f_reg(370) <= "00010101000101100000000000110101";
                        f_reg(371) <= "10101111101010000000011111100100";
                        f_reg(372) <= "10001100000111010000100001000000";
                        f_reg(373) <= "00011111101000000000000000000011";
                        f_reg(374) <= "00100000000111010000000000111100";
                        f_reg(375) <= "00010000000000000000000000000010";
                        f_reg(376) <= "00100000000111010000000000000000";
                        f_reg(377) <= "00010101001101110000000000101110";
                        f_reg(378) <= "10101111101010010000011111101000";
                        f_reg(379) <= "10001100000111010000100001000000";
                        f_reg(380) <= "00011111101000000000000000000011";
                        f_reg(381) <= "00100000000111010000000000111100";
                        f_reg(382) <= "00010000000000000000000000000010";
                        f_reg(383) <= "00100000000111010000000000000000";
                        f_reg(384) <= "00010101010110000000000000100111";
                        f_reg(385) <= "10101111101010100000011111101100";
                        f_reg(386) <= "10001100000111010000100001000000";
                        f_reg(387) <= "00011111101000000000000000000011";
                        f_reg(388) <= "00100000000111010000000000111100";
                        f_reg(389) <= "00010000000000000000000000000010";
                        f_reg(390) <= "00100000000111010000000000000000";
                        f_reg(391) <= "00010101011110010000000000100000";
                        f_reg(392) <= "10101111101010110000011111110000";
                        f_reg(393) <= "10001100000111010000100001000000";
                        f_reg(394) <= "00011111101000000000000000000011";
                        f_reg(395) <= "00100000000111010000000000111100";
                        f_reg(396) <= "00010000000000000000000000000010";
                        f_reg(397) <= "00100000000111010000000000000000";
                        f_reg(398) <= "00010101100110100000000000011001";
                        f_reg(399) <= "10101111101011000000011111110100";
                        f_reg(400) <= "10001100000111010000100001000000";
                        f_reg(401) <= "00011111101000000000000000000011";
                        f_reg(402) <= "00100000000111010000000000111100";
                        f_reg(403) <= "00010000000000000000000000000010";
                        f_reg(404) <= "00100000000111010000000000000000";
                        f_reg(405) <= "00010101101110110000000000010010";
                        f_reg(406) <= "10101111101011010000011111111000";
                        f_reg(407) <= "10001100000111010000100001000000";
                        f_reg(408) <= "00011111101000000000000000000011";
                        f_reg(409) <= "00100000000111010000000000111100";
                        f_reg(410) <= "00010000000000000000000000000010";
                        f_reg(411) <= "00100000000111010000000000000000";
                        f_reg(412) <= "00010101110111000000000000001011";
                        f_reg(413) <= "10101111101011100000011111111100";
                        f_reg(414) <= "10001100000111010000100001000000";
                        f_reg(415) <= "00011111101000000000000000000011";
                        f_reg(416) <= "00100000000111010000000000111100";
                        f_reg(417) <= "00010000000000000000000000000010";
                        f_reg(418) <= "00100000000111010000000000000000";
                        f_reg(419) <= "00010111110111110000000000000100";
                        f_reg(420) <= "10101111101111100000100000000000";
                        f_reg(421) <= "10101100000111010000100001000000";
                        f_reg(422) <= "00010000000000001111111101111011";
                        f_reg(423) <= "10001100000111010000100001000000";
                        f_reg(424) <= "10001111101000010000011111001000";
                        f_reg(425) <= "10001100000111010000100001000000";
                        f_reg(426) <= "10001111101011110000011111001000";
                        f_reg(427) <= "00010100001011111111111111111100";
                        f_reg(428) <= "10001100000111010000100001000000";
                        f_reg(429) <= "10001111101000100000011111001100";
                        f_reg(430) <= "10001100000111010000100001000000";
                        f_reg(431) <= "10001111101100000000011111001100";
                        f_reg(432) <= "00010100010100001111111111111100";
                        f_reg(433) <= "10001100000111010000100001000000";
                        f_reg(434) <= "10001111101000110000011111010000";
                        f_reg(435) <= "10001100000111010000100001000000";
                        f_reg(436) <= "10001111101100010000011111010000";
                        f_reg(437) <= "00010100011100011111111111111100";
                        f_reg(438) <= "10001100000111010000100001000000";
                        f_reg(439) <= "10001111101001000000011111010100";
                        f_reg(440) <= "10001100000111010000100001000000";
                        f_reg(441) <= "10001111101100100000011111010100";
                        f_reg(442) <= "00010100100100101111111111111100";
                        f_reg(443) <= "10001100000111010000100001000000";
                        f_reg(444) <= "10001111101001010000011111011000";
                        f_reg(445) <= "10001100000111010000100001000000";
                        f_reg(446) <= "10001111101100110000011111011000";
                        f_reg(447) <= "00010100101100111111111111111100";
                        f_reg(448) <= "10001100000111010000100001000000";
                        f_reg(449) <= "10001111101001100000011111011100";
                        f_reg(450) <= "10001100000111010000100001000000";
                        f_reg(451) <= "10001111101101000000011111011100";
                        f_reg(452) <= "00010100110101001111111111111100";
                        f_reg(453) <= "10001100000111010000100001000000";
                        f_reg(454) <= "10001111101001110000011111100000";
                        f_reg(455) <= "10001100000111010000100001000000";
                        f_reg(456) <= "10001111101101010000011111100000";
                        f_reg(457) <= "00010100111101011111111111111100";
                        f_reg(458) <= "10001100000111010000100001000000";
                        f_reg(459) <= "10001111101010000000011111100100";
                        f_reg(460) <= "10001100000111010000100001000000";
                        f_reg(461) <= "10001111101101100000011111100100";
                        f_reg(462) <= "00010101000101101111111111111100";
                        f_reg(463) <= "10001100000111010000100001000000";
                        f_reg(464) <= "10001111101010010000011111101000";
                        f_reg(465) <= "10001100000111010000100001000000";
                        f_reg(466) <= "10001111101101110000011111101000";
                        f_reg(467) <= "00010101001101111111111111111100";
                        f_reg(468) <= "10001100000111010000100001000000";
                        f_reg(469) <= "10001111101010100000011111101100";
                        f_reg(470) <= "10001100000111010000100001000000";
                        f_reg(471) <= "10001111101110000000011111101100";
                        f_reg(472) <= "00010101010110001111111111111100";
                        f_reg(473) <= "10001100000111010000100001000000";
                        f_reg(474) <= "10001111101010110000011111110000";
                        f_reg(475) <= "10001100000111010000100001000000";
                        f_reg(476) <= "10001111101110010000011111110000";
                        f_reg(477) <= "00010101011110011111111111111100";
                        f_reg(478) <= "10001100000111010000100001000000";
                        f_reg(479) <= "10001111101011000000011111110100";
                        f_reg(480) <= "10001100000111010000100001000000";
                        f_reg(481) <= "10001111101110100000011111110100";
                        f_reg(482) <= "00010101100110101111111111111100";
                        f_reg(483) <= "10001100000111010000100001000000";
                        f_reg(484) <= "10001111101011010000011111111000";
                        f_reg(485) <= "10001100000111010000100001000000";
                        f_reg(486) <= "10001111101110110000011111111000";
                        f_reg(487) <= "00010101101110111111111111111100";
                        f_reg(488) <= "10001100000111010000100001000000";
                        f_reg(489) <= "10001111101011100000011111111100";
                        f_reg(490) <= "10001100000111010000100001000000";
                        f_reg(491) <= "10001111101111000000011111111100";
                        f_reg(492) <= "00010101110111001111111111111100";
                        f_reg(493) <= "10001100000111010000100001000000";
                        f_reg(494) <= "10001111101111100000100000000000";
                        f_reg(495) <= "10001100000111010000100001000000";
                        f_reg(496) <= "10001111101111110000100000000000";
                        f_reg(497) <= "00010111110111111111111111111100";
                        f_reg(498) <= "00010000000000001111111100101111";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000001111100111";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                        f_reg(551) <= "00000000000000000000000000000000";
                        f_reg(552) <= "00000000000000000000000000000000";
                        f_reg(553) <= "00000000000000000000000000000000";
                        f_reg(554) <= "00000000000000000000000000000000";
                        f_reg(555) <= "00000000000000000000000000000000";
                        f_reg(556) <= "00000000000000000000000000000000";
                        f_reg(557) <= "00000000000000000000000000000000";
                        f_reg(558) <= "00000000000000000000000000000000";
                        f_reg(559) <= "00000000000000000000000000000000";
                        f_reg(560) <= "00000000000000000000000000000000";
                        f_reg(561) <= "00000000000000000000000000000000";
                        f_reg(562) <= "00000000000000000000000000000000";
                        f_reg(563) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 3914
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- XORI R2 R0 -13506
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- SW R1 R0 1172
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SRL R3 R0 20
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SUBU R4 R1 R2
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- XORI R5 R2 11459
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- ANDI R6 R4 23545
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- ADD R7 R2 R6
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- SUB R8 R3 R2
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- ADDIU R9 R4 -9117
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- ANDI R10 R3 7716
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- SRLV R11 R8 R8
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- SW R6 R0 1176
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- ADD R12 R6 R9
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- ADD R13 R9 R8
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- SRLV R14 R12 R1
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SRLV R15 R10 R14
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- SLTI R16 R11 11687
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- SW R1 R0 1180
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- SRLV R17 R4 R9
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- SLLV R18 R7 R1
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- SW R6 R0 1184
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- NOP
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- SRL R19 R12 5
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- SUB R20 R18 R6
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- NOR R21 R11 R16
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- SW R13 R0 1188
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- AND R22 R16 R9
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- OR R23 R4 R18
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- XOR R24 R17 R19
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- LUI R25 2845
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- SUB R26 R25 R19
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- SRL R27 R17 2
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- SLLV R28 R26 R26
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- NOR R29 R0 R28
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- SLTIU R30 R24 -30200
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- NOR R2 R22 R20
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- ADDU R3 R27 R15
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- LUI R8 14691
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- NOR R14 R30 R25
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SRL R7 R10 14
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- ADD R6 R22 R0
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- NOP
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- ADDIU R13 R25 -2004
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- SLTI R16 R30 7583
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- ADD R9 R26 R21
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- ADDU R4 R11 R23
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- OR R18 R13 R9
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- SRAV R19 R8 R7
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- ADDU R17 R2 R3
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- NOP
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SLTIU R1 R1 6520
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SW R6 R0 1192
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- AND R24 R18 R5
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SW R24 R0 1196
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- ADD R27 R28 R16
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- ADD R15 R27 R21
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- SRA R10 R21 27
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- SLLV R10 R10 R4
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- SLT R22 R20 R12
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- SLTU R25 R29 R17
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- SW R21 R0 1200
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- ANDI R30 R10 -23233
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- SRLV R26 R14 R19
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- NOR R11 R25 R22
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- ADDI R23 R11 -10409
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- SLTI R13 R30 7371
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SW R26 R0 1204
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- SW R22 R0 1208
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- SW R15 R0 1212
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SW R26 R0 1216
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- XORI R9 R25 -16469
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- SLTI R8 R23 -20018
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- SW R1 R0 1220
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- SW R8 R0 1224
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- ADDI R7 R9 13692
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- SW R19 R0 1228
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- AND R2 R7 R23
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- ADDI R3 R2 4706
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- SW R13 R0 1232
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SW R3 R0 1236
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- ADDI R31 R31 -1
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- BGTZ R31 -82
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- BEQ R0 R0 478
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- LUI R30 999
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- LUI R31 999
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- SRL R30 R30 16
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- SRL R31 R31 16
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- LUI R1 3914
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- LUI R15 3914
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- XORI R2 R0 -13506
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- XORI R16 R0 -13506
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- BNE R1 R15 328
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- SW R1 R0 1172
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SRL R3 R0 20
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SRL R17 R0 20
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- SUBU R4 R1 R2
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- SUBU R18 R15 R16
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- XORI R5 R2 11459
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- XORI R19 R16 11459
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- ANDI R6 R4 23545
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- ANDI R20 R18 23545
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- ADD R7 R2 R6
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- ADD R21 R16 R20
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- SUB R8 R3 R2
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- SUB R22 R17 R16
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- ADDIU R9 R4 -9117
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- ADDIU R23 R18 -9117
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- ANDI R10 R3 7716
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- ANDI R24 R17 7716
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- SRLV R11 R8 R8
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- SRLV R25 R22 R22
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- BNE R6 R20 308
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- SW R6 R0 1176
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- ADD R12 R6 R9
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- ADD R26 R20 R23
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- ADD R13 R9 R8
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- ADD R27 R23 R22
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- SRLV R14 R12 R1
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- SRLV R28 R26 R15
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- SRLV R2 R10 R14
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SRLV R16 R24 R28
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- SLTI R3 R11 11687
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- SLTI R17 R25 11687
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- BNE R1 R15 296
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SW R1 R0 1180
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- SRLV R8 R4 R9
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- SRLV R22 R18 R23
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- SLLV R14 R7 R1
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- SLLV R28 R21 R15
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- BNE R6 R20 290
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- SW R6 R0 1184
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- NOP
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- NOP
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- SRL R7 R12 5
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SRL R21 R26 5
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- BNE R12 R26 284
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- SW R12 R0 1240
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- SUB R12 R14 R6
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- SUB R26 R28 R20
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- NOR R6 R11 R3
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- NOR R20 R25 R17
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- BNE R13 R27 278
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- SW R13 R0 1188
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- AND R13 R3 R9
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- AND R27 R17 R23
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- OR R3 R4 R14
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- OR R17 R18 R28
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- XOR R9 R8 R7
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- XOR R23 R22 R21
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- LUI R4 2845
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- LUI R18 2845
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- SUB R14 R4 R7
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- SUB R28 R18 R21
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- SRL R7 R8 2
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- SRL R21 R22 2
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- SLLV R8 R14 R14
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- SLLV R22 R28 R28
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- BNE R6 R20 262
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- SW R6 R0 1244
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- NOR R6 R0 R8
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- NOR R20 R0 R22
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- BNE R6 R20 258
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- SW R6 R0 1248
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- SLTIU R6 R9 -30200
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- SLTIU R20 R23 -30200
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- NOR R9 R13 R12
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- NOR R23 R27 R26
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- BNE R12 R26 252
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- SW R12 R0 1252
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- ADDU R12 R7 R2
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- ADDU R26 R21 R16
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- LUI R7 14691
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- LUI R21 14691
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- NOR R2 R6 R4
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- NOR R16 R20 R18
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- BNE R2 R16 244
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- SW R2 R0 1256
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- SRL R2 R10 14
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SRL R16 R24 14
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- ADD R10 R13 R0
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- ADD R24 R27 R0
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- NOP
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- NOP
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- ADDIU R13 R4 -2004
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- ADDIU R27 R18 -2004
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- SLTI R4 R6 7583
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- SLTI R18 R20 7583
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- LW R6 R0 1244
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- LW R20 R0 1244
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- BNE R6 R20 -2
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- BNE R8 R22 229
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- SW R8 R0 1244
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- ADD R8 R14 R6
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- ADD R22 R28 R20
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- ADDU R14 R11 R3
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- ADDU R28 R25 R17
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- OR R11 R13 R8
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- OR R25 R27 R22
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- SRAV R3 R7 R2
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- SRAV R17 R21 R16
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- ADDU R13 R9 R12
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- ADDU R27 R23 R26
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- NOP
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- NOP
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- SLTIU R1 R1 6520
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- SLTIU R15 R15 6520
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- BNE R10 R24 213
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- SW R10 R0 1192
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- AND R8 R11 R5
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- AND R22 R25 R19
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- BNE R8 R22 209
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- SW R8 R0 1196
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- LW R7 R0 1244
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- LW R21 R0 1244
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- BNE R7 R21 -2
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- ADD R2 R7 R4
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- ADD R16 R21 R18
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- ADD R9 R2 R6
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- ADD R23 R16 R20
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- SRA R12 R6 27
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- SRA R26 R20 27
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- SLLV R12 R12 R14
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- SLLV R26 R26 R28
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- LW R10 R0 1252
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- LW R24 R0 1252
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- BNE R10 R24 -2
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- LW R11 R0 1240
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- LW R25 R0 1240
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- BNE R11 R25 -2
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- SLT R5 R10 R11
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- SLT R19 R24 R25
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- LW R8 R0 1248
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- LW R22 R0 1248
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- BNE R8 R22 -2
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- SLTU R7 R8 R13
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- SLTU R21 R22 R27
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- BNE R6 R20 183
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- SW R6 R0 1200
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- ANDI R4 R12 -23233
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- ANDI R18 R26 -23233
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- LW R2 R0 1256
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- LW R16 R0 1256
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- BNE R2 R16 -2
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- SRLV R14 R2 R3
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- SRLV R28 R16 R17
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- NOR R10 R7 R5
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- NOR R24 R21 R19
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- ADDI R11 R10 -10409
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- ADDI R25 R24 -10409
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- SLTI R8 R4 7371
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- SLTI R22 R18 7371
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- BNE R14 R28 168
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- SW R14 R0 1204
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- BNE R5 R19 166
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- SW R5 R0 1208
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- BNE R9 R23 164
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- SW R9 R0 1212
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- BNE R14 R28 162
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- SW R14 R0 1216
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- XORI R13 R7 -16469
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- XORI R27 R21 -16469
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- SLTI R6 R11 -20018
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- SLTI R20 R25 -20018
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- BNE R1 R15 156
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- SW R1 R0 1220
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- BNE R6 R20 154
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- SW R6 R0 1224
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- ADDI R12 R13 13692
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- ADDI R26 R27 13692
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- BNE R3 R17 150
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- SW R3 R0 1228
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- AND R2 R12 R11
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- AND R16 R26 R25
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- ADDI R10 R2 4706
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- ADDI R24 R16 4706
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- BNE R8 R22 144
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- SW R8 R0 1232
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- BNE R10 R24 142
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- SW R10 R0 1236
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- ADDI R29 R30 -250
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- BEQ R29 R0 32
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- ADDI R29 R30 -500
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- BEQ R29 R0 30
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- ADDI R29 R30 -750
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- BEQ R29 R0 28
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- ADDI R30 R30 -1
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- ADDI R31 R31 -1
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- BNE R30 R31 132
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- BGTZ R31 -201
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- BEQ R0 R0 271
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- NOP
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- NOP
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- NOP
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- NOP
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- NOP
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- NOP
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- NOP
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- NOP
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- NOP
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- NOP
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- NOP
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- NOP
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- NOP
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- NOP
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- NOP
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- NOP
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- NOP
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- NOP
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- NOP
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- NOP
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- NOP
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- NOP
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- LW R29 R0 2112
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- BGTZ R29 3
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- ADDI R29 R0 60
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- BEQ R0 R0 2
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- ADDI R29 R0 0
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- BNE R1 R15 102
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- SW R1 R29 1992
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- LW R29 R0 2112
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- BGTZ R29 3
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- ADDI R29 R0 60
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- BEQ R0 R0 2
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- ADDI R29 R0 0
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- BNE R2 R16 95
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- SW R2 R29 1996
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- LW R29 R0 2112
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- BGTZ R29 3
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- ADDI R29 R0 60
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- BEQ R0 R0 2
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- ADDI R29 R0 0
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- BNE R3 R17 88
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- SW R3 R29 2000
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- LW R29 R0 2112
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- BGTZ R29 3
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- ADDI R29 R0 60
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- BEQ R0 R0 2
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- ADDI R29 R0 0
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- BNE R4 R18 81
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- SW R4 R29 2004
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- LW R29 R0 2112
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- BGTZ R29 3
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- ADDI R29 R0 60
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- BEQ R0 R0 2
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- ADDI R29 R0 0
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- BNE R5 R19 74
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- SW R5 R29 2008
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- LW R29 R0 2112
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- BGTZ R29 3
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- ADDI R29 R0 60
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- BEQ R0 R0 2
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- ADDI R29 R0 0
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- BNE R6 R20 67
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- SW R6 R29 2012
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- LW R29 R0 2112
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- BGTZ R29 3
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- ADDI R29 R0 60
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- BEQ R0 R0 2
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- ADDI R29 R0 0
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- BNE R7 R21 60
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- SW R7 R29 2016
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- LW R29 R0 2112
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- BGTZ R29 3
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- ADDI R29 R0 60
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- BEQ R0 R0 2
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- ADDI R29 R0 0
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- BNE R8 R22 53
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- SW R8 R29 2020
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- LW R29 R0 2112
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- BGTZ R29 3
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- ADDI R29 R0 60
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- BEQ R0 R0 2
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- ADDI R29 R0 0
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- BNE R9 R23 46
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- SW R9 R29 2024
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- LW R29 R0 2112
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- BGTZ R29 3
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- ADDI R29 R0 60
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- BEQ R0 R0 2
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- ADDI R29 R0 0
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- BNE R10 R24 39
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- SW R10 R29 2028
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- LW R29 R0 2112
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- BGTZ R29 3
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- ADDI R29 R0 60
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- BEQ R0 R0 2
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- ADDI R29 R0 0
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- BNE R11 R25 32
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- SW R11 R29 2032
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- LW R29 R0 2112
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- BGTZ R29 3
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- ADDI R29 R0 60
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- BEQ R0 R0 2
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- ADDI R29 R0 0
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- BNE R12 R26 25
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- SW R12 R29 2036
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- LW R29 R0 2112
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- BGTZ R29 3
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- ADDI R29 R0 60
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- BEQ R0 R0 2
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- ADDI R29 R0 0
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- BNE R13 R27 18
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- SW R13 R29 2040
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- LW R29 R0 2112
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- BGTZ R29 3
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- ADDI R29 R0 60
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- BEQ R0 R0 2
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- ADDI R29 R0 0
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- BNE R14 R28 11
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- SW R14 R29 2044
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- LW R29 R0 2112
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- BGTZ R29 3
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- ADDI R29 R0 60
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- BEQ R0 R0 2
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- ADDI R29 R0 0
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- BNE R30 R31 4
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- SW R30 R29 2048
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- SW R29 R0 2112
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- BEQ R0 R0 -133
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- LW R29 R0 2112
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- LW R1 R29 1992
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R29 R0 2112
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R15 R29 1992
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- BNE R1 R15 -4
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- LW R29 R0 2112
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- LW R2 R29 1996
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- LW R29 R0 2112
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- LW R16 R29 1996
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- BNE R2 R16 -4
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- LW R29 R0 2112
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- LW R3 R29 2000
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- LW R29 R0 2112
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- LW R17 R29 2000
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- BNE R3 R17 -4
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- LW R29 R0 2112
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- LW R4 R29 2004
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- LW R29 R0 2112
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- LW R18 R29 2004
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- BNE R4 R18 -4
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- LW R29 R0 2112
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- LW R5 R29 2008
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- LW R29 R0 2112
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- LW R19 R29 2008
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- BNE R5 R19 -4
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- LW R29 R0 2112
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- LW R6 R29 2012
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- LW R29 R0 2112
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- LW R20 R29 2012
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- BNE R6 R20 -4
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- LW R29 R0 2112
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- LW R7 R29 2016
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- LW R29 R0 2112
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- LW R21 R29 2016
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- BNE R7 R21 -4
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- LW R29 R0 2112
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- LW R8 R29 2020
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- LW R29 R0 2112
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- LW R22 R29 2020
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- BNE R8 R22 -4
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- LW R29 R0 2112
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- LW R9 R29 2024
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- LW R29 R0 2112
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- LW R23 R29 2024
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- BNE R9 R23 -4
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- LW R29 R0 2112
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- LW R10 R29 2028
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- LW R29 R0 2112
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- LW R24 R29 2028
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- BNE R10 R24 -4
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- LW R29 R0 2112
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- LW R11 R29 2032
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- LW R29 R0 2112
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- LW R25 R29 2032
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- BNE R11 R25 -4
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- LW R29 R0 2112
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- LW R12 R29 2036
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- LW R29 R0 2112
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- LW R26 R29 2036
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- BNE R12 R26 -4
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- LW R29 R0 2112
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- LW R13 R29 2040
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- LW R29 R0 2112
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- LW R27 R29 2040
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- BNE R13 R27 -4
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- LW R29 R0 2112
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- LW R14 R29 2044
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- LW R29 R0 2112
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- LW R28 R29 2044
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- BNE R14 R28 -4
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- LW R29 R0 2112
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- LW R30 R29 2048
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- LW R29 R0 2112
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- LW R31 R29 2048
                        f_reg(496) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(497) =>
                        -- BNE R30 R31 -4
                        f_reg(497) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(498) =>
                        -- BEQ R0 R0 -209
                        f_reg(498) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(499) =>
                        -- NOP
                        f_reg(499) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(500) =>
                        -- NOP
                        f_reg(500) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(501) =>
                        -- NOP
                        f_reg(501) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(502) =>
                        -- NOP
                        f_reg(502) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(503) =>
                        -- NOP
                        f_reg(503) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(504) =>
                        -- NOP
                        f_reg(504) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(505) =>
                        -- NOP
                        f_reg(505) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(506) =>
                        -- NOP
                        f_reg(506) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(507) =>
                        -- NOP
                        f_reg(507) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(508) =>
                        -- NOP
                        f_reg(508) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(509) =>
                        -- NOP
                        f_reg(509) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(510) =>
                        -- NOP
                        f_reg(510) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(511) =>
                        -- NOP
                        f_reg(511) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(512) =>
                        -- NOP
                        f_reg(512) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(513) =>
                        -- NOP
                        f_reg(513) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(514) =>
                        -- NOP
                        f_reg(514) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(515) =>
                        -- NOP
                        f_reg(515) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(516) =>
                        -- NOP
                        f_reg(516) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(517) =>
                        -- NOP
                        f_reg(517) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(518) =>
                        -- NOP
                        f_reg(518) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(519) =>
                        -- NOP
                        f_reg(519) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(520) =>
                        -- NOP
                        f_reg(520) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(521) =>
                        -- NOP
                        f_reg(521) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(522) =>
                        -- NOP
                        f_reg(522) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(523) =>
                        -- NOP
                        f_reg(523) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(524) =>
                        -- NOP
                        f_reg(524) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(525) =>
                        -- NOP
                        f_reg(525) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(526) =>
                        -- NOP
                        f_reg(526) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(527) =>
                        -- NOP
                        f_reg(527) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(528) =>
                        -- NOP
                        f_reg(528) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(529) =>
                        -- NOP
                        f_reg(529) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(530) =>
                        -- NOP
                        f_reg(530) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(531) =>
                        -- NOP
                        f_reg(531) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(532) =>
                        -- NOP
                        f_reg(532) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(533) =>
                        -- NOP
                        f_reg(533) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(534) =>
                        -- NOP
                        f_reg(534) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(535) =>
                        -- NOP
                        f_reg(535) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(536) =>
                        -- NOP
                        f_reg(536) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(537) =>
                        -- NOP
                        f_reg(537) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(538) =>
                        -- NOP
                        f_reg(538) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(539) =>
                        -- NOP
                        f_reg(539) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(540) =>
                        -- NOP
                        f_reg(540) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(541) =>
                        -- NOP
                        f_reg(541) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(542) =>
                        -- NOP
                        f_reg(542) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(543) =>
                        -- NOP
                        f_reg(543) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(544) =>
                        -- NOP
                        f_reg(544) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(545) =>
                        -- NOP
                        f_reg(545) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(546) =>
                        -- NOP
                        f_reg(546) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(547) =>
                        -- NOP
                        f_reg(547) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(548) =>
                        -- NOP
                        f_reg(548) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(549) =>
                        -- NOP
                        f_reg(549) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(550) =>
                        -- NOP
                        f_reg(550) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(551) =>
                        -- NOP
                        f_reg(551) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(552) =>
                        -- NOP
                        f_reg(552) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(553) =>
                        -- NOP
                        f_reg(553) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(554) =>
                        -- NOP
                        f_reg(554) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(555) =>
                        -- NOP
                        f_reg(555) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(556) =>
                        -- NOP
                        f_reg(556) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(557) =>
                        -- NOP
                        f_reg(557) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(558) =>
                        -- NOP
                        f_reg(558) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(559) =>
                        -- NOP
                        f_reg(559) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(560) =>
                        -- NOP
                        f_reg(560) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(561) =>
                        -- NOP
                        f_reg(561) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(562) =>
                        -- NOP
                        f_reg(562) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(563) =>
                        -- NOP
                        f_reg(563) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(564) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010000111101001010";
                        f_reg(4) <= "00111000000000101100101100111110";
                        f_reg(5) <= "10101100000000010000010010010100";
                        f_reg(6) <= "00000000000000000001110100000010";
                        f_reg(7) <= "00000000001000100010000000100011";
                        f_reg(8) <= "00111000010001010010110011000011";
                        f_reg(9) <= "00110000100001100101101111111001";
                        f_reg(10) <= "00000000010001100011100000100000";
                        f_reg(11) <= "00000000011000100100000000100010";
                        f_reg(12) <= "00100100100010011101110001100011";
                        f_reg(13) <= "00110000011010100001111000100100";
                        f_reg(14) <= "00000001000010000101100000000110";
                        f_reg(15) <= "10101100000001100000010010011000";
                        f_reg(16) <= "00000000110010010110000000100000";
                        f_reg(17) <= "00000001001010000110100000100000";
                        f_reg(18) <= "00000000001011000111000000000110";
                        f_reg(19) <= "00000001110010100111100000000110";
                        f_reg(20) <= "00101001011100000010110110100111";
                        f_reg(21) <= "10101100000000010000010010011100";
                        f_reg(22) <= "00000001001001001000100000000110";
                        f_reg(23) <= "00000000001001111001000000000100";
                        f_reg(24) <= "10101100000001100000010010100000";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00000000000011001001100101000010";
                        f_reg(27) <= "00000010010001101010000000100010";
                        f_reg(28) <= "00000001011100001010100000100111";
                        f_reg(29) <= "10101100000011010000010010100100";
                        f_reg(30) <= "00000010000010011011000000100100";
                        f_reg(31) <= "00000000100100101011100000100101";
                        f_reg(32) <= "00000010001100111100000000100110";
                        f_reg(33) <= "00111100000110010000101100011101";
                        f_reg(34) <= "00000011001100111101000000100010";
                        f_reg(35) <= "00000000000100011101100010000010";
                        f_reg(36) <= "00000011010110101110000000000100";
                        f_reg(37) <= "00000000000111001110100000100111";
                        f_reg(38) <= "00101111000111101000101000001000";
                        f_reg(39) <= "00000010110101000001000000100111";
                        f_reg(40) <= "00000011011011110001100000100001";
                        f_reg(41) <= "00111100000010000011100101100011";
                        f_reg(42) <= "00000011110110010111000000100111";
                        f_reg(43) <= "00000000000010100011101110000010";
                        f_reg(44) <= "00000010110000000011000000100000";
                        f_reg(45) <= "00000000000000000000000000000000";
                        f_reg(46) <= "00100111001011011111100000101100";
                        f_reg(47) <= "00101011110100000001110110011111";
                        f_reg(48) <= "00000011010101010100100000100000";
                        f_reg(49) <= "00000001011101110010000000100001";
                        f_reg(50) <= "00000001101010011001000000100101";
                        f_reg(51) <= "00000000111010001001100000000111";
                        f_reg(52) <= "00000000010000111000100000100001";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00101100001000010001100101111000";
                        f_reg(55) <= "10101100000001100000010010101000";
                        f_reg(56) <= "00000010010001011100000000100100";
                        f_reg(57) <= "10101100000110000000010010101100";
                        f_reg(58) <= "00000011100100001101100000100000";
                        f_reg(59) <= "00000011011101010111100000100000";
                        f_reg(60) <= "00000000000101010101011011000011";
                        f_reg(61) <= "00000000100010100101000000000100";
                        f_reg(62) <= "00000010100011001011000000101010";
                        f_reg(63) <= "00000011101100011100100000101011";
                        f_reg(64) <= "10101100000101010000010010110000";
                        f_reg(65) <= "00110001010111101010010100111111";
                        f_reg(66) <= "00000010011011101101000000000110";
                        f_reg(67) <= "00000011001101100101100000100111";
                        f_reg(68) <= "00100001011101111101011101010111";
                        f_reg(69) <= "00101011110011010001110011001011";
                        f_reg(70) <= "10101100000110100000010010110100";
                        f_reg(71) <= "10101100000101100000010010111000";
                        f_reg(72) <= "10101100000011110000010010111100";
                        f_reg(73) <= "10101100000110100000010011000000";
                        f_reg(74) <= "00111011001010011011111110101011";
                        f_reg(75) <= "00101010111010001011000111001110";
                        f_reg(76) <= "10101100000000010000010011000100";
                        f_reg(77) <= "10101100000010000000010011001000";
                        f_reg(78) <= "00100001001001110011010101111100";
                        f_reg(79) <= "10101100000100110000010011001100";
                        f_reg(80) <= "00000000111101110001000000100100";
                        f_reg(81) <= "00100000010000110001001001100010";
                        f_reg(82) <= "10101100000011010000010011010000";
                        f_reg(83) <= "10101100000000110000010011010100";
                        f_reg(84) <= "00100011111111111111111111111111";
                        f_reg(85) <= "00011111111000001111111110101110";
                        f_reg(86) <= "00010000000000000000000111011110";
                        f_reg(87) <= "00111100000111100000001111100111";
                        f_reg(88) <= "00111100000111110000001111100111";
                        f_reg(89) <= "00000000000111101111010000000010";
                        f_reg(90) <= "00000000000111111111110000000010";
                        f_reg(91) <= "00111100000000010000111101001010";
                        f_reg(92) <= "00111100000011110000111101001010";
                        f_reg(93) <= "00111000000000101100101100111110";
                        f_reg(94) <= "00111000000100001100101100111110";
                        f_reg(95) <= "00010100001011110000000101001000";
                        f_reg(96) <= "10101100000000010000010010010100";
                        f_reg(97) <= "00000000000000000001110100000010";
                        f_reg(98) <= "00000000000000001000110100000010";
                        f_reg(99) <= "00000000001000100010000000100011";
                        f_reg(100) <= "00000001111100001001000000100011";
                        f_reg(101) <= "00111000010001010010110011000011";
                        f_reg(102) <= "00111010000100110010110011000011";
                        f_reg(103) <= "00110000100001100101101111111001";
                        f_reg(104) <= "00110010010101000101101111111001";
                        f_reg(105) <= "00000000010001100011100000100000";
                        f_reg(106) <= "00000010000101001010100000100000";
                        f_reg(107) <= "00000000011000100100000000100010";
                        f_reg(108) <= "00000010001100001011000000100010";
                        f_reg(109) <= "00100100100010011101110001100011";
                        f_reg(110) <= "00100110010101111101110001100011";
                        f_reg(111) <= "00110000011010100001111000100100";
                        f_reg(112) <= "00110010001110000001111000100100";
                        f_reg(113) <= "00000001000010000101100000000110";
                        f_reg(114) <= "00000010110101101100100000000110";
                        f_reg(115) <= "00010100110101000000000100110100";
                        f_reg(116) <= "10101100000001100000010010011000";
                        f_reg(117) <= "00000000110010010110000000100000";
                        f_reg(118) <= "00000010100101111101000000100000";
                        f_reg(119) <= "00000001001010000110100000100000";
                        f_reg(120) <= "00000010111101101101100000100000";
                        f_reg(121) <= "00000000001011000111000000000110";
                        f_reg(122) <= "00000001111110101110000000000110";
                        f_reg(123) <= "00000001110010100001000000000110";
                        f_reg(124) <= "00000011100110001000000000000110";
                        f_reg(125) <= "00101001011000110010110110100111";
                        f_reg(126) <= "00101011001100010010110110100111";
                        f_reg(127) <= "00010100001011110000000100101000";
                        f_reg(128) <= "10101100000000010000010010011100";
                        f_reg(129) <= "00000001001001000100000000000110";
                        f_reg(130) <= "00000010111100101011000000000110";
                        f_reg(131) <= "00000000001001110111000000000100";
                        f_reg(132) <= "00000001111101011110000000000100";
                        f_reg(133) <= "00010100110101000000000100100010";
                        f_reg(134) <= "10101100000001100000010010100000";
                        f_reg(135) <= "00000000000000000000000000000000";
                        f_reg(136) <= "00000000000000000000000000000000";
                        f_reg(137) <= "00000000000011000011100101000010";
                        f_reg(138) <= "00000000000110101010100101000010";
                        f_reg(139) <= "00010101100110100000000100011100";
                        f_reg(140) <= "10101100000011000000010011011000";
                        f_reg(141) <= "00000001110001100110000000100010";
                        f_reg(142) <= "00000011100101001101000000100010";
                        f_reg(143) <= "00000001011000110011000000100111";
                        f_reg(144) <= "00000011001100011010000000100111";
                        f_reg(145) <= "00010101101110110000000100010110";
                        f_reg(146) <= "10101100000011010000010010100100";
                        f_reg(147) <= "00000000011010010110100000100100";
                        f_reg(148) <= "00000010001101111101100000100100";
                        f_reg(149) <= "00000000100011100001100000100101";
                        f_reg(150) <= "00000010010111001000100000100101";
                        f_reg(151) <= "00000001000001110100100000100110";
                        f_reg(152) <= "00000010110101011011100000100110";
                        f_reg(153) <= "00111100000001000000101100011101";
                        f_reg(154) <= "00111100000100100000101100011101";
                        f_reg(155) <= "00000000100001110111000000100010";
                        f_reg(156) <= "00000010010101011110000000100010";
                        f_reg(157) <= "00000000000010000011100010000010";
                        f_reg(158) <= "00000000000101101010100010000010";
                        f_reg(159) <= "00000001110011100100000000000100";
                        f_reg(160) <= "00000011100111001011000000000100";
                        f_reg(161) <= "00010100110101000000000100000110";
                        f_reg(162) <= "10101100000001100000010011011100";
                        f_reg(163) <= "00000000000010000011000000100111";
                        f_reg(164) <= "00000000000101101010000000100111";
                        f_reg(165) <= "00010100110101000000000100000010";
                        f_reg(166) <= "10101100000001100000010011100000";
                        f_reg(167) <= "00101101001001101000101000001000";
                        f_reg(168) <= "00101110111101001000101000001000";
                        f_reg(169) <= "00000001101011000100100000100111";
                        f_reg(170) <= "00000011011110101011100000100111";
                        f_reg(171) <= "00010101100110100000000011111100";
                        f_reg(172) <= "10101100000011000000010011100100";
                        f_reg(173) <= "00000000111000100110000000100001";
                        f_reg(174) <= "00000010101100001101000000100001";
                        f_reg(175) <= "00111100000001110011100101100011";
                        f_reg(176) <= "00111100000101010011100101100011";
                        f_reg(177) <= "00000000110001000001000000100111";
                        f_reg(178) <= "00000010100100101000000000100111";
                        f_reg(179) <= "00010100010100000000000011110100";
                        f_reg(180) <= "10101100000000100000010011101000";
                        f_reg(181) <= "00000000000010100001001110000010";
                        f_reg(182) <= "00000000000110001000001110000010";
                        f_reg(183) <= "00000001101000000101000000100000";
                        f_reg(184) <= "00000011011000001100000000100000";
                        f_reg(185) <= "00000000000000000000000000000000";
                        f_reg(186) <= "00000000000000000000000000000000";
                        f_reg(187) <= "00100100100011011111100000101100";
                        f_reg(188) <= "00100110010110111111100000101100";
                        f_reg(189) <= "00101000110001000001110110011111";
                        f_reg(190) <= "00101010100100100001110110011111";
                        f_reg(191) <= "10001100000001100000010011011100";
                        f_reg(192) <= "10001100000101000000010011011100";
                        f_reg(193) <= "00010100110101001111111111111110";
                        f_reg(194) <= "00010101000101100000000011100101";
                        f_reg(195) <= "10101100000010000000010011011100";
                        f_reg(196) <= "00000001110001100100000000100000";
                        f_reg(197) <= "00000011100101001011000000100000";
                        f_reg(198) <= "00000001011000110111000000100001";
                        f_reg(199) <= "00000011001100011110000000100001";
                        f_reg(200) <= "00000001101010000101100000100101";
                        f_reg(201) <= "00000011011101101100100000100101";
                        f_reg(202) <= "00000000010001110001100000000111";
                        f_reg(203) <= "00000010000101011000100000000111";
                        f_reg(204) <= "00000001001011000110100000100001";
                        f_reg(205) <= "00000010111110101101100000100001";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101100001000010001100101111000";
                        f_reg(209) <= "00101101111011110001100101111000";
                        f_reg(210) <= "00010101010110000000000011010101";
                        f_reg(211) <= "10101100000010100000010010101000";
                        f_reg(212) <= "00000001011001010100000000100100";
                        f_reg(213) <= "00000011001100111011000000100100";
                        f_reg(214) <= "00010101000101100000000011010001";
                        f_reg(215) <= "10101100000010000000010010101100";
                        f_reg(216) <= "10001100000001110000010011011100";
                        f_reg(217) <= "10001100000101010000010011011100";
                        f_reg(218) <= "00010100111101011111111111111110";
                        f_reg(219) <= "00000000111001000001000000100000";
                        f_reg(220) <= "00000010101100101000000000100000";
                        f_reg(221) <= "00000000010001100100100000100000";
                        f_reg(222) <= "00000010000101001011100000100000";
                        f_reg(223) <= "00000000000001100110011011000011";
                        f_reg(224) <= "00000000000101001101011011000011";
                        f_reg(225) <= "00000001110011000110000000000100";
                        f_reg(226) <= "00000011100110101101000000000100";
                        f_reg(227) <= "10001100000010100000010011100100";
                        f_reg(228) <= "10001100000110000000010011100100";
                        f_reg(229) <= "00010101010110001111111111111110";
                        f_reg(230) <= "10001100000010110000010011011000";
                        f_reg(231) <= "10001100000110010000010011011000";
                        f_reg(232) <= "00010101011110011111111111111110";
                        f_reg(233) <= "00000001010010110010100000101010";
                        f_reg(234) <= "00000011000110011001100000101010";
                        f_reg(235) <= "10001100000010000000010011100000";
                        f_reg(236) <= "10001100000101100000010011100000";
                        f_reg(237) <= "00010101000101101111111111111110";
                        f_reg(238) <= "00000001000011010011100000101011";
                        f_reg(239) <= "00000010110110111010100000101011";
                        f_reg(240) <= "00010100110101000000000010110111";
                        f_reg(241) <= "10101100000001100000010010110000";
                        f_reg(242) <= "00110001100001001010010100111111";
                        f_reg(243) <= "00110011010100101010010100111111";
                        f_reg(244) <= "10001100000000100000010011101000";
                        f_reg(245) <= "10001100000100000000010011101000";
                        f_reg(246) <= "00010100010100001111111111111110";
                        f_reg(247) <= "00000000011000100111000000000110";
                        f_reg(248) <= "00000010001100001110000000000110";
                        f_reg(249) <= "00000000111001010101000000100111";
                        f_reg(250) <= "00000010101100111100000000100111";
                        f_reg(251) <= "00100001010010111101011101010111";
                        f_reg(252) <= "00100011000110011101011101010111";
                        f_reg(253) <= "00101000100010000001110011001011";
                        f_reg(254) <= "00101010010101100001110011001011";
                        f_reg(255) <= "00010101110111000000000010101000";
                        f_reg(256) <= "10101100000011100000010010110100";
                        f_reg(257) <= "00010100101100110000000010100110";
                        f_reg(258) <= "10101100000001010000010010111000";
                        f_reg(259) <= "00010101001101110000000010100100";
                        f_reg(260) <= "10101100000010010000010010111100";
                        f_reg(261) <= "00010101110111000000000010100010";
                        f_reg(262) <= "10101100000011100000010011000000";
                        f_reg(263) <= "00111000111011011011111110101011";
                        f_reg(264) <= "00111010101110111011111110101011";
                        f_reg(265) <= "00101001011001101011000111001110";
                        f_reg(266) <= "00101011001101001011000111001110";
                        f_reg(267) <= "00010100001011110000000010011100";
                        f_reg(268) <= "10101100000000010000010011000100";
                        f_reg(269) <= "00010100110101000000000010011010";
                        f_reg(270) <= "10101100000001100000010011001000";
                        f_reg(271) <= "00100001101011000011010101111100";
                        f_reg(272) <= "00100011011110100011010101111100";
                        f_reg(273) <= "00010100011100010000000010010110";
                        f_reg(274) <= "10101100000000110000010011001100";
                        f_reg(275) <= "00000001100010110001000000100100";
                        f_reg(276) <= "00000011010110011000000000100100";
                        f_reg(277) <= "00100000010010100001001001100010";
                        f_reg(278) <= "00100010000110000001001001100010";
                        f_reg(279) <= "00010101000101100000000010010000";
                        f_reg(280) <= "10101100000010000000010011010000";
                        f_reg(281) <= "00010101010110000000000010001110";
                        f_reg(282) <= "10101100000010100000010011010100";
                        f_reg(283) <= "00100011110111011111111100000110";
                        f_reg(284) <= "00010011101000000000000000100000";
                        f_reg(285) <= "00100011110111011111111000001100";
                        f_reg(286) <= "00010011101000000000000000011110";
                        f_reg(287) <= "00100011110111011111110100010010";
                        f_reg(288) <= "00010011101000000000000000011100";
                        f_reg(289) <= "00100011110111101111111111111111";
                        f_reg(290) <= "00100011111111111111111111111111";
                        f_reg(291) <= "00010111110111110000000010000100";
                        f_reg(292) <= "00011111111000001111111100110111";
                        f_reg(293) <= "00010000000000000000000100001111";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "00000000000000000000000000000000";
                        f_reg(304) <= "00000000000000000000000000000000";
                        f_reg(305) <= "00000000000000000000000000000000";
                        f_reg(306) <= "00000000000000000000000000000000";
                        f_reg(307) <= "00000000000000000000000000000000";
                        f_reg(308) <= "00000000000000000000000000000000";
                        f_reg(309) <= "00000000000000000000000000000000";
                        f_reg(310) <= "00000000000000000000000000000000";
                        f_reg(311) <= "00000000000000000000000000000000";
                        f_reg(312) <= "00000000000000000000000000000000";
                        f_reg(313) <= "00000000000000000000000000000000";
                        f_reg(314) <= "00000000000000000000000000000000";
                        f_reg(315) <= "00000000000000000000000000000000";
                        f_reg(316) <= "10001100000111010000100001000000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010100001011110000000001100110";
                        f_reg(322) <= "10101111101000010000011111001000";
                        f_reg(323) <= "10001100000111010000100001000000";
                        f_reg(324) <= "00011111101000000000000000000011";
                        f_reg(325) <= "00100000000111010000000000111100";
                        f_reg(326) <= "00010000000000000000000000000010";
                        f_reg(327) <= "00100000000111010000000000000000";
                        f_reg(328) <= "00010100010100000000000001011111";
                        f_reg(329) <= "10101111101000100000011111001100";
                        f_reg(330) <= "10001100000111010000100001000000";
                        f_reg(331) <= "00011111101000000000000000000011";
                        f_reg(332) <= "00100000000111010000000000111100";
                        f_reg(333) <= "00010000000000000000000000000010";
                        f_reg(334) <= "00100000000111010000000000000000";
                        f_reg(335) <= "00010100011100010000000001011000";
                        f_reg(336) <= "10101111101000110000011111010000";
                        f_reg(337) <= "10001100000111010000100001000000";
                        f_reg(338) <= "00011111101000000000000000000011";
                        f_reg(339) <= "00100000000111010000000000111100";
                        f_reg(340) <= "00010000000000000000000000000010";
                        f_reg(341) <= "00100000000111010000000000000000";
                        f_reg(342) <= "00010100100100100000000001010001";
                        f_reg(343) <= "10101111101001000000011111010100";
                        f_reg(344) <= "10001100000111010000100001000000";
                        f_reg(345) <= "00011111101000000000000000000011";
                        f_reg(346) <= "00100000000111010000000000111100";
                        f_reg(347) <= "00010000000000000000000000000010";
                        f_reg(348) <= "00100000000111010000000000000000";
                        f_reg(349) <= "00010100101100110000000001001010";
                        f_reg(350) <= "10101111101001010000011111011000";
                        f_reg(351) <= "10001100000111010000100001000000";
                        f_reg(352) <= "00011111101000000000000000000011";
                        f_reg(353) <= "00100000000111010000000000111100";
                        f_reg(354) <= "00010000000000000000000000000010";
                        f_reg(355) <= "00100000000111010000000000000000";
                        f_reg(356) <= "00010100110101000000000001000011";
                        f_reg(357) <= "10101111101001100000011111011100";
                        f_reg(358) <= "10001100000111010000100001000000";
                        f_reg(359) <= "00011111101000000000000000000011";
                        f_reg(360) <= "00100000000111010000000000111100";
                        f_reg(361) <= "00010000000000000000000000000010";
                        f_reg(362) <= "00100000000111010000000000000000";
                        f_reg(363) <= "00010100111101010000000000111100";
                        f_reg(364) <= "10101111101001110000011111100000";
                        f_reg(365) <= "10001100000111010000100001000000";
                        f_reg(366) <= "00011111101000000000000000000011";
                        f_reg(367) <= "00100000000111010000000000111100";
                        f_reg(368) <= "00010000000000000000000000000010";
                        f_reg(369) <= "00100000000111010000000000000000";
                        f_reg(370) <= "00010101000101100000000000110101";
                        f_reg(371) <= "10101111101010000000011111100100";
                        f_reg(372) <= "10001100000111010000100001000000";
                        f_reg(373) <= "00011111101000000000000000000011";
                        f_reg(374) <= "00100000000111010000000000111100";
                        f_reg(375) <= "00010000000000000000000000000010";
                        f_reg(376) <= "00100000000111010000000000000000";
                        f_reg(377) <= "00010101001101110000000000101110";
                        f_reg(378) <= "10101111101010010000011111101000";
                        f_reg(379) <= "10001100000111010000100001000000";
                        f_reg(380) <= "00011111101000000000000000000011";
                        f_reg(381) <= "00100000000111010000000000111100";
                        f_reg(382) <= "00010000000000000000000000000010";
                        f_reg(383) <= "00100000000111010000000000000000";
                        f_reg(384) <= "00010101010110000000000000100111";
                        f_reg(385) <= "10101111101010100000011111101100";
                        f_reg(386) <= "10001100000111010000100001000000";
                        f_reg(387) <= "00011111101000000000000000000011";
                        f_reg(388) <= "00100000000111010000000000111100";
                        f_reg(389) <= "00010000000000000000000000000010";
                        f_reg(390) <= "00100000000111010000000000000000";
                        f_reg(391) <= "00010101011110010000000000100000";
                        f_reg(392) <= "10101111101010110000011111110000";
                        f_reg(393) <= "10001100000111010000100001000000";
                        f_reg(394) <= "00011111101000000000000000000011";
                        f_reg(395) <= "00100000000111010000000000111100";
                        f_reg(396) <= "00010000000000000000000000000010";
                        f_reg(397) <= "00100000000111010000000000000000";
                        f_reg(398) <= "00010101100110100000000000011001";
                        f_reg(399) <= "10101111101011000000011111110100";
                        f_reg(400) <= "10001100000111010000100001000000";
                        f_reg(401) <= "00011111101000000000000000000011";
                        f_reg(402) <= "00100000000111010000000000111100";
                        f_reg(403) <= "00010000000000000000000000000010";
                        f_reg(404) <= "00100000000111010000000000000000";
                        f_reg(405) <= "00010101101110110000000000010010";
                        f_reg(406) <= "10101111101011010000011111111000";
                        f_reg(407) <= "10001100000111010000100001000000";
                        f_reg(408) <= "00011111101000000000000000000011";
                        f_reg(409) <= "00100000000111010000000000111100";
                        f_reg(410) <= "00010000000000000000000000000010";
                        f_reg(411) <= "00100000000111010000000000000000";
                        f_reg(412) <= "00010101110111000000000000001011";
                        f_reg(413) <= "10101111101011100000011111111100";
                        f_reg(414) <= "10001100000111010000100001000000";
                        f_reg(415) <= "00011111101000000000000000000011";
                        f_reg(416) <= "00100000000111010000000000111100";
                        f_reg(417) <= "00010000000000000000000000000010";
                        f_reg(418) <= "00100000000111010000000000000000";
                        f_reg(419) <= "00010111110111110000000000000100";
                        f_reg(420) <= "10101111101111100000100000000000";
                        f_reg(421) <= "10101100000111010000100001000000";
                        f_reg(422) <= "00010000000000001111111101111011";
                        f_reg(423) <= "10001100000111010000100001000000";
                        f_reg(424) <= "10001111101000010000011111001000";
                        f_reg(425) <= "10001100000111010000100001000000";
                        f_reg(426) <= "10001111101011110000011111001000";
                        f_reg(427) <= "00010100001011111111111111111100";
                        f_reg(428) <= "10001100000111010000100001000000";
                        f_reg(429) <= "10001111101000100000011111001100";
                        f_reg(430) <= "10001100000111010000100001000000";
                        f_reg(431) <= "10001111101100000000011111001100";
                        f_reg(432) <= "00010100010100001111111111111100";
                        f_reg(433) <= "10001100000111010000100001000000";
                        f_reg(434) <= "10001111101000110000011111010000";
                        f_reg(435) <= "10001100000111010000100001000000";
                        f_reg(436) <= "10001111101100010000011111010000";
                        f_reg(437) <= "00010100011100011111111111111100";
                        f_reg(438) <= "10001100000111010000100001000000";
                        f_reg(439) <= "10001111101001000000011111010100";
                        f_reg(440) <= "10001100000111010000100001000000";
                        f_reg(441) <= "10001111101100100000011111010100";
                        f_reg(442) <= "00010100100100101111111111111100";
                        f_reg(443) <= "10001100000111010000100001000000";
                        f_reg(444) <= "10001111101001010000011111011000";
                        f_reg(445) <= "10001100000111010000100001000000";
                        f_reg(446) <= "10001111101100110000011111011000";
                        f_reg(447) <= "00010100101100111111111111111100";
                        f_reg(448) <= "10001100000111010000100001000000";
                        f_reg(449) <= "10001111101001100000011111011100";
                        f_reg(450) <= "10001100000111010000100001000000";
                        f_reg(451) <= "10001111101101000000011111011100";
                        f_reg(452) <= "00010100110101001111111111111100";
                        f_reg(453) <= "10001100000111010000100001000000";
                        f_reg(454) <= "10001111101001110000011111100000";
                        f_reg(455) <= "10001100000111010000100001000000";
                        f_reg(456) <= "10001111101101010000011111100000";
                        f_reg(457) <= "00010100111101011111111111111100";
                        f_reg(458) <= "10001100000111010000100001000000";
                        f_reg(459) <= "10001111101010000000011111100100";
                        f_reg(460) <= "10001100000111010000100001000000";
                        f_reg(461) <= "10001111101101100000011111100100";
                        f_reg(462) <= "00010101000101101111111111111100";
                        f_reg(463) <= "10001100000111010000100001000000";
                        f_reg(464) <= "10001111101010010000011111101000";
                        f_reg(465) <= "10001100000111010000100001000000";
                        f_reg(466) <= "10001111101101110000011111101000";
                        f_reg(467) <= "00010101001101111111111111111100";
                        f_reg(468) <= "10001100000111010000100001000000";
                        f_reg(469) <= "10001111101010100000011111101100";
                        f_reg(470) <= "10001100000111010000100001000000";
                        f_reg(471) <= "10001111101110000000011111101100";
                        f_reg(472) <= "00010101010110001111111111111100";
                        f_reg(473) <= "10001100000111010000100001000000";
                        f_reg(474) <= "10001111101010110000011111110000";
                        f_reg(475) <= "10001100000111010000100001000000";
                        f_reg(476) <= "10001111101110010000011111110000";
                        f_reg(477) <= "00010101011110011111111111111100";
                        f_reg(478) <= "10001100000111010000100001000000";
                        f_reg(479) <= "10001111101011000000011111110100";
                        f_reg(480) <= "10001100000111010000100001000000";
                        f_reg(481) <= "10001111101110100000011111110100";
                        f_reg(482) <= "00010101100110101111111111111100";
                        f_reg(483) <= "10001100000111010000100001000000";
                        f_reg(484) <= "10001111101011010000011111111000";
                        f_reg(485) <= "10001100000111010000100001000000";
                        f_reg(486) <= "10001111101110110000011111111000";
                        f_reg(487) <= "00010101101110111111111111111100";
                        f_reg(488) <= "10001100000111010000100001000000";
                        f_reg(489) <= "10001111101011100000011111111100";
                        f_reg(490) <= "10001100000111010000100001000000";
                        f_reg(491) <= "10001111101111000000011111111100";
                        f_reg(492) <= "00010101110111001111111111111100";
                        f_reg(493) <= "10001100000111010000100001000000";
                        f_reg(494) <= "10001111101111100000100000000000";
                        f_reg(495) <= "10001100000111010000100001000000";
                        f_reg(496) <= "10001111101111110000100000000000";
                        f_reg(497) <= "00010111110111111111111111111100";
                        f_reg(498) <= "00010000000000001111111100101111";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000001111100111";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                        f_reg(551) <= "00000000000000000000000000000000";
                        f_reg(552) <= "00000000000000000000000000000000";
                        f_reg(553) <= "00000000000000000000000000000000";
                        f_reg(554) <= "00000000000000000000000000000000";
                        f_reg(555) <= "00000000000000000000000000000000";
                        f_reg(556) <= "00000000000000000000000000000000";
                        f_reg(557) <= "00000000000000000000000000000000";
                        f_reg(558) <= "00000000000000000000000000000000";
                        f_reg(559) <= "00000000000000000000000000000000";
                        f_reg(560) <= "00000000000000000000000000000000";
                        f_reg(561) <= "00000000000000000000000000000000";
                        f_reg(562) <= "00000000000000000000000000000000";
                        f_reg(563) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000010000111101001010";
                        f_reg(4) <= "00111000000000101100101100111110";
                        f_reg(5) <= "10101100000000010000010010010100";
                        f_reg(6) <= "00000000000000000001110100000010";
                        f_reg(7) <= "00000000001000100010000000100011";
                        f_reg(8) <= "00111000010001010010110011000011";
                        f_reg(9) <= "00110000100001100101101111111001";
                        f_reg(10) <= "00000000010001100011100000100000";
                        f_reg(11) <= "00000000011000100100000000100010";
                        f_reg(12) <= "00100100100010011101110001100011";
                        f_reg(13) <= "00110000011010100001111000100100";
                        f_reg(14) <= "00000001000010000101100000000110";
                        f_reg(15) <= "10101100000001100000010010011000";
                        f_reg(16) <= "00000000110010010110000000100000";
                        f_reg(17) <= "00000001001010000110100000100000";
                        f_reg(18) <= "00000000001011000111000000000110";
                        f_reg(19) <= "00000001110010100111100000000110";
                        f_reg(20) <= "00101001011100000010110110100111";
                        f_reg(21) <= "10101100000000010000010010011100";
                        f_reg(22) <= "00000001001001001000100000000110";
                        f_reg(23) <= "00000000001001111001000000000100";
                        f_reg(24) <= "10101100000001100000010010100000";
                        f_reg(25) <= "00000000000000000000000000000000";
                        f_reg(26) <= "00000000000011001001100101000010";
                        f_reg(27) <= "00000010010001101010000000100010";
                        f_reg(28) <= "00000001011100001010100000100111";
                        f_reg(29) <= "10101100000011010000010010100100";
                        f_reg(30) <= "00000010000010011011000000100100";
                        f_reg(31) <= "00000000100100101011100000100101";
                        f_reg(32) <= "00000010001100111100000000100110";
                        f_reg(33) <= "00111100000110010000101100011101";
                        f_reg(34) <= "00000011001100111101000000100010";
                        f_reg(35) <= "00000000000100011101100010000010";
                        f_reg(36) <= "00000011010110101110000000000100";
                        f_reg(37) <= "00000000000111001110100000100111";
                        f_reg(38) <= "00101111000111101000101000001000";
                        f_reg(39) <= "00000010110101000001000000100111";
                        f_reg(40) <= "00000011011011110001100000100001";
                        f_reg(41) <= "00111100000010000011100101100011";
                        f_reg(42) <= "00000011110110010111000000100111";
                        f_reg(43) <= "00000000000010100011101110000010";
                        f_reg(44) <= "00000010110000000011000000100000";
                        f_reg(45) <= "00000000000000000000000000000000";
                        f_reg(46) <= "00100111001011011111100000101100";
                        f_reg(47) <= "00101011110100000001110110011111";
                        f_reg(48) <= "00000011010101010100100000100000";
                        f_reg(49) <= "00000001011101110010000000100001";
                        f_reg(50) <= "00000001101010011001000000100101";
                        f_reg(51) <= "00000000111010001001100000000111";
                        f_reg(52) <= "00000000010000111000100000100001";
                        f_reg(53) <= "00000000000000000000000000000000";
                        f_reg(54) <= "00101100001000010001100101111000";
                        f_reg(55) <= "10101100000001100000010010101000";
                        f_reg(56) <= "00000010010001011100000000100100";
                        f_reg(57) <= "10101100000110000000010010101100";
                        f_reg(58) <= "00000011100100001101100000100000";
                        f_reg(59) <= "00000011011101010111100000100000";
                        f_reg(60) <= "00000000000101010101011011000011";
                        f_reg(61) <= "00000000100010100101000000000100";
                        f_reg(62) <= "00000010100011001011000000101010";
                        f_reg(63) <= "00000011101100011100100000101011";
                        f_reg(64) <= "10101100000101010000010010110000";
                        f_reg(65) <= "00110001010111101010010100111111";
                        f_reg(66) <= "00000010011011101101000000000110";
                        f_reg(67) <= "00000011001101100101100000100111";
                        f_reg(68) <= "00100001011101111101011101010111";
                        f_reg(69) <= "00101011110011010001110011001011";
                        f_reg(70) <= "10101100000110100000010010110100";
                        f_reg(71) <= "10101100000101100000010010111000";
                        f_reg(72) <= "10101100000011110000010010111100";
                        f_reg(73) <= "10101100000110100000010011000000";
                        f_reg(74) <= "00111011001010011011111110101011";
                        f_reg(75) <= "00101010111010001011000111001110";
                        f_reg(76) <= "10101100000000010000010011000100";
                        f_reg(77) <= "10101100000010000000010011001000";
                        f_reg(78) <= "00100001001001110011010101111100";
                        f_reg(79) <= "10101100000100110000010011001100";
                        f_reg(80) <= "00000000111101110001000000100100";
                        f_reg(81) <= "00100000010000110001001001100010";
                        f_reg(82) <= "10101100000011010000010011010000";
                        f_reg(83) <= "10101100000000110000010011010100";
                        f_reg(84) <= "00100011111111111111111111111111";
                        f_reg(85) <= "00011111111000001111111110101110";
                        f_reg(86) <= "00010000000000000000000111011110";
                        f_reg(87) <= "00111100000111100000001111100111";
                        f_reg(88) <= "00111100000111110000001111100111";
                        f_reg(89) <= "00000000000111101111010000000010";
                        f_reg(90) <= "00000000000111111111110000000010";
                        f_reg(91) <= "00111100000000010000111101001010";
                        f_reg(92) <= "00111100000011110000111101001010";
                        f_reg(93) <= "00111000000000101100101100111110";
                        f_reg(94) <= "00111000000100001100101100111110";
                        f_reg(95) <= "00010100001011110000000101001000";
                        f_reg(96) <= "10101100000000010000010010010100";
                        f_reg(97) <= "00000000000000000001110100000010";
                        f_reg(98) <= "00000000000000001000110100000010";
                        f_reg(99) <= "00000000001000100010000000100011";
                        f_reg(100) <= "00000001111100001001000000100011";
                        f_reg(101) <= "00111000010001010010110011000011";
                        f_reg(102) <= "00111010000100110010110011000011";
                        f_reg(103) <= "00110000100001100101101111111001";
                        f_reg(104) <= "00110010010101000101101111111001";
                        f_reg(105) <= "00000000010001100011100000100000";
                        f_reg(106) <= "00000010000101001010100000100000";
                        f_reg(107) <= "00000000011000100100000000100010";
                        f_reg(108) <= "00000010001100001011000000100010";
                        f_reg(109) <= "00100100100010011101110001100011";
                        f_reg(110) <= "00100110010101111101110001100011";
                        f_reg(111) <= "00110000011010100001111000100100";
                        f_reg(112) <= "00110010001110000001111000100100";
                        f_reg(113) <= "00000001000010000101100000000110";
                        f_reg(114) <= "00000010110101101100100000000110";
                        f_reg(115) <= "00010100110101000000000100110100";
                        f_reg(116) <= "10101100000001100000010010011000";
                        f_reg(117) <= "00000000110010010110000000100000";
                        f_reg(118) <= "00000010100101111101000000100000";
                        f_reg(119) <= "00000001001010000110100000100000";
                        f_reg(120) <= "00000010111101101101100000100000";
                        f_reg(121) <= "00000000001011000111000000000110";
                        f_reg(122) <= "00000001111110101110000000000110";
                        f_reg(123) <= "00000001110010100001000000000110";
                        f_reg(124) <= "00000011100110001000000000000110";
                        f_reg(125) <= "00101001011000110010110110100111";
                        f_reg(126) <= "00101011001100010010110110100111";
                        f_reg(127) <= "00010100001011110000000100101000";
                        f_reg(128) <= "10101100000000010000010010011100";
                        f_reg(129) <= "00000001001001000100000000000110";
                        f_reg(130) <= "00000010111100101011000000000110";
                        f_reg(131) <= "00000000001001110111000000000100";
                        f_reg(132) <= "00000001111101011110000000000100";
                        f_reg(133) <= "00010100110101000000000100100010";
                        f_reg(134) <= "10101100000001100000010010100000";
                        f_reg(135) <= "00000000000000000000000000000000";
                        f_reg(136) <= "00000000000000000000000000000000";
                        f_reg(137) <= "00000000000011000011100101000010";
                        f_reg(138) <= "00000000000110101010100101000010";
                        f_reg(139) <= "00010101100110100000000100011100";
                        f_reg(140) <= "10101100000011000000010011011000";
                        f_reg(141) <= "00000001110001100110000000100010";
                        f_reg(142) <= "00000011100101001101000000100010";
                        f_reg(143) <= "00000001011000110011000000100111";
                        f_reg(144) <= "00000011001100011010000000100111";
                        f_reg(145) <= "00010101101110110000000100010110";
                        f_reg(146) <= "10101100000011010000010010100100";
                        f_reg(147) <= "00000000011010010110100000100100";
                        f_reg(148) <= "00000010001101111101100000100100";
                        f_reg(149) <= "00000000100011100001100000100101";
                        f_reg(150) <= "00000010010111001000100000100101";
                        f_reg(151) <= "00000001000001110100100000100110";
                        f_reg(152) <= "00000010110101011011100000100110";
                        f_reg(153) <= "00111100000001000000101100011101";
                        f_reg(154) <= "00111100000100100000101100011101";
                        f_reg(155) <= "00000000100001110111000000100010";
                        f_reg(156) <= "00000010010101011110000000100010";
                        f_reg(157) <= "00000000000010000011100010000010";
                        f_reg(158) <= "00000000000101101010100010000010";
                        f_reg(159) <= "00000001110011100100000000000100";
                        f_reg(160) <= "00000011100111001011000000000100";
                        f_reg(161) <= "00010100110101000000000100000110";
                        f_reg(162) <= "10101100000001100000010011011100";
                        f_reg(163) <= "00000000000010000011000000100111";
                        f_reg(164) <= "00000000000101101010000000100111";
                        f_reg(165) <= "00010100110101000000000100000010";
                        f_reg(166) <= "10101100000001100000010011100000";
                        f_reg(167) <= "00101101001001101000101000001000";
                        f_reg(168) <= "00101110111101001000101000001000";
                        f_reg(169) <= "00000001101011000100100000100111";
                        f_reg(170) <= "00000011011110101011100000100111";
                        f_reg(171) <= "00010101100110100000000011111100";
                        f_reg(172) <= "10101100000011000000010011100100";
                        f_reg(173) <= "00000000111000100110000000100001";
                        f_reg(174) <= "00000010101100001101000000100001";
                        f_reg(175) <= "00111100000001110011100101100011";
                        f_reg(176) <= "00111100000101010011100101100011";
                        f_reg(177) <= "00000000110001000001000000100111";
                        f_reg(178) <= "00000010100100101000000000100111";
                        f_reg(179) <= "00010100010100000000000011110100";
                        f_reg(180) <= "10101100000000100000010011101000";
                        f_reg(181) <= "00000000000010100001001110000010";
                        f_reg(182) <= "00000000000110001000001110000010";
                        f_reg(183) <= "00000001101000000101000000100000";
                        f_reg(184) <= "00000011011000001100000000100000";
                        f_reg(185) <= "00000000000000000000000000000000";
                        f_reg(186) <= "00000000000000000000000000000000";
                        f_reg(187) <= "00100100100011011111100000101100";
                        f_reg(188) <= "00100110010110111111100000101100";
                        f_reg(189) <= "00101000110001000001110110011111";
                        f_reg(190) <= "00101010100100100001110110011111";
                        f_reg(191) <= "10001100000001100000010011011100";
                        f_reg(192) <= "10001100000101000000010011011100";
                        f_reg(193) <= "00010100110101001111111111111110";
                        f_reg(194) <= "00010101000101100000000011100101";
                        f_reg(195) <= "10101100000010000000010011011100";
                        f_reg(196) <= "00000001110001100100000000100000";
                        f_reg(197) <= "00000011100101001011000000100000";
                        f_reg(198) <= "00000001011000110111000000100001";
                        f_reg(199) <= "00000011001100011110000000100001";
                        f_reg(200) <= "00000001101010000101100000100101";
                        f_reg(201) <= "00000011011101101100100000100101";
                        f_reg(202) <= "00000000010001110001100000000111";
                        f_reg(203) <= "00000010000101011000100000000111";
                        f_reg(204) <= "00000001001011000110100000100001";
                        f_reg(205) <= "00000010111110101101100000100001";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101100001000010001100101111000";
                        f_reg(209) <= "00101101111011110001100101111000";
                        f_reg(210) <= "00010101010110000000000011010101";
                        f_reg(211) <= "10101100000010100000010010101000";
                        f_reg(212) <= "00000001011001010100000000100100";
                        f_reg(213) <= "00000011001100111011000000100100";
                        f_reg(214) <= "00010101000101100000000011010001";
                        f_reg(215) <= "10101100000010000000010010101100";
                        f_reg(216) <= "10001100000001110000010011011100";
                        f_reg(217) <= "10001100000101010000010011011100";
                        f_reg(218) <= "00010100111101011111111111111110";
                        f_reg(219) <= "00000000111001000001000000100000";
                        f_reg(220) <= "00000010101100101000000000100000";
                        f_reg(221) <= "00000000010001100100100000100000";
                        f_reg(222) <= "00000010000101001011100000100000";
                        f_reg(223) <= "00000000000001100110011011000011";
                        f_reg(224) <= "00000000000101001101011011000011";
                        f_reg(225) <= "00000001110011000110000000000100";
                        f_reg(226) <= "00000011100110101101000000000100";
                        f_reg(227) <= "10001100000010100000010011100100";
                        f_reg(228) <= "10001100000110000000010011100100";
                        f_reg(229) <= "00010101010110001111111111111110";
                        f_reg(230) <= "10001100000010110000010011011000";
                        f_reg(231) <= "10001100000110010000010011011000";
                        f_reg(232) <= "00010101011110011111111111111110";
                        f_reg(233) <= "00000001010010110010100000101010";
                        f_reg(234) <= "00000011000110011001100000101010";
                        f_reg(235) <= "10001100000010000000010011100000";
                        f_reg(236) <= "10001100000101100000010011100000";
                        f_reg(237) <= "00010101000101101111111111111110";
                        f_reg(238) <= "00000001000011010011100000101011";
                        f_reg(239) <= "00000010110110111010100000101011";
                        f_reg(240) <= "00010100110101000000000010110111";
                        f_reg(241) <= "10101100000001100000010010110000";
                        f_reg(242) <= "00110001100001001010010100111111";
                        f_reg(243) <= "00110011010100101010010100111111";
                        f_reg(244) <= "10001100000000100000010011101000";
                        f_reg(245) <= "10001100000100000000010011101000";
                        f_reg(246) <= "00010100010100001111111111111110";
                        f_reg(247) <= "00000000011000100111000000000110";
                        f_reg(248) <= "00000010001100001110000000000110";
                        f_reg(249) <= "00000000111001010101000000100111";
                        f_reg(250) <= "00000010101100111100000000100111";
                        f_reg(251) <= "00100001010010111101011101010111";
                        f_reg(252) <= "00100011000110011101011101010111";
                        f_reg(253) <= "00101000100010000001110011001011";
                        f_reg(254) <= "00101010010101100001110011001011";
                        f_reg(255) <= "00010101110111000000000010101000";
                        f_reg(256) <= "10101100000011100000010010110100";
                        f_reg(257) <= "00010100101100110000000010100110";
                        f_reg(258) <= "10101100000001010000010010111000";
                        f_reg(259) <= "00010101001101110000000010100100";
                        f_reg(260) <= "10101100000010010000010010111100";
                        f_reg(261) <= "00010101110111000000000010100010";
                        f_reg(262) <= "10101100000011100000010011000000";
                        f_reg(263) <= "00111000111011011011111110101011";
                        f_reg(264) <= "00111010101110111011111110101011";
                        f_reg(265) <= "00101001011001101011000111001110";
                        f_reg(266) <= "00101011001101001011000111001110";
                        f_reg(267) <= "00010100001011110000000010011100";
                        f_reg(268) <= "10101100000000010000010011000100";
                        f_reg(269) <= "00010100110101000000000010011010";
                        f_reg(270) <= "10101100000001100000010011001000";
                        f_reg(271) <= "00100001101011000011010101111100";
                        f_reg(272) <= "00100011011110100011010101111100";
                        f_reg(273) <= "00010100011100010000000010010110";
                        f_reg(274) <= "10101100000000110000010011001100";
                        f_reg(275) <= "00000001100010110001000000100100";
                        f_reg(276) <= "00000011010110011000000000100100";
                        f_reg(277) <= "00100000010010100001001001100010";
                        f_reg(278) <= "00100010000110000001001001100010";
                        f_reg(279) <= "00010101000101100000000010010000";
                        f_reg(280) <= "10101100000010000000010011010000";
                        f_reg(281) <= "00010101010110000000000010001110";
                        f_reg(282) <= "10101100000010100000010011010100";
                        f_reg(283) <= "00100011110111011111111100000110";
                        f_reg(284) <= "00010011101000000000000000100000";
                        f_reg(285) <= "00100011110111011111111000001100";
                        f_reg(286) <= "00010011101000000000000000011110";
                        f_reg(287) <= "00100011110111011111110100010010";
                        f_reg(288) <= "00010011101000000000000000011100";
                        f_reg(289) <= "00100011110111101111111111111111";
                        f_reg(290) <= "00100011111111111111111111111111";
                        f_reg(291) <= "00010111110111110000000010000100";
                        f_reg(292) <= "00011111111000001111111100110111";
                        f_reg(293) <= "00010000000000000000000100001111";
                        f_reg(294) <= "00000000000000000000000000000000";
                        f_reg(295) <= "00000000000000000000000000000000";
                        f_reg(296) <= "00000000000000000000000000000000";
                        f_reg(297) <= "00000000000000000000000000000000";
                        f_reg(298) <= "00000000000000000000000000000000";
                        f_reg(299) <= "00000000000000000000000000000000";
                        f_reg(300) <= "00000000000000000000000000000000";
                        f_reg(301) <= "00000000000000000000000000000000";
                        f_reg(302) <= "00000000000000000000000000000000";
                        f_reg(303) <= "00000000000000000000000000000000";
                        f_reg(304) <= "00000000000000000000000000000000";
                        f_reg(305) <= "00000000000000000000000000000000";
                        f_reg(306) <= "00000000000000000000000000000000";
                        f_reg(307) <= "00000000000000000000000000000000";
                        f_reg(308) <= "00000000000000000000000000000000";
                        f_reg(309) <= "00000000000000000000000000000000";
                        f_reg(310) <= "00000000000000000000000000000000";
                        f_reg(311) <= "00000000000000000000000000000000";
                        f_reg(312) <= "00000000000000000000000000000000";
                        f_reg(313) <= "00000000000000000000000000000000";
                        f_reg(314) <= "00000000000000000000000000000000";
                        f_reg(315) <= "00000000000000000000000000000000";
                        f_reg(316) <= "10001100000111010000100001000000";
                        f_reg(317) <= "00011111101000000000000000000011";
                        f_reg(318) <= "00100000000111010000000000111100";
                        f_reg(319) <= "00010000000000000000000000000010";
                        f_reg(320) <= "00100000000111010000000000000000";
                        f_reg(321) <= "00010100001011110000000001100110";
                        f_reg(322) <= "10101111101000010000011111001000";
                        f_reg(323) <= "10001100000111010000100001000000";
                        f_reg(324) <= "00011111101000000000000000000011";
                        f_reg(325) <= "00100000000111010000000000111100";
                        f_reg(326) <= "00010000000000000000000000000010";
                        f_reg(327) <= "00100000000111010000000000000000";
                        f_reg(328) <= "00010100010100000000000001011111";
                        f_reg(329) <= "10101111101000100000011111001100";
                        f_reg(330) <= "10001100000111010000100001000000";
                        f_reg(331) <= "00011111101000000000000000000011";
                        f_reg(332) <= "00100000000111010000000000111100";
                        f_reg(333) <= "00010000000000000000000000000010";
                        f_reg(334) <= "00100000000111010000000000000000";
                        f_reg(335) <= "00010100011100010000000001011000";
                        f_reg(336) <= "10101111101000110000011111010000";
                        f_reg(337) <= "10001100000111010000100001000000";
                        f_reg(338) <= "00011111101000000000000000000011";
                        f_reg(339) <= "00100000000111010000000000111100";
                        f_reg(340) <= "00010000000000000000000000000010";
                        f_reg(341) <= "00100000000111010000000000000000";
                        f_reg(342) <= "00010100100100100000000001010001";
                        f_reg(343) <= "10101111101001000000011111010100";
                        f_reg(344) <= "10001100000111010000100001000000";
                        f_reg(345) <= "00011111101000000000000000000011";
                        f_reg(346) <= "00100000000111010000000000111100";
                        f_reg(347) <= "00010000000000000000000000000010";
                        f_reg(348) <= "00100000000111010000000000000000";
                        f_reg(349) <= "00010100101100110000000001001010";
                        f_reg(350) <= "10101111101001010000011111011000";
                        f_reg(351) <= "10001100000111010000100001000000";
                        f_reg(352) <= "00011111101000000000000000000011";
                        f_reg(353) <= "00100000000111010000000000111100";
                        f_reg(354) <= "00010000000000000000000000000010";
                        f_reg(355) <= "00100000000111010000000000000000";
                        f_reg(356) <= "00010100110101000000000001000011";
                        f_reg(357) <= "10101111101001100000011111011100";
                        f_reg(358) <= "10001100000111010000100001000000";
                        f_reg(359) <= "00011111101000000000000000000011";
                        f_reg(360) <= "00100000000111010000000000111100";
                        f_reg(361) <= "00010000000000000000000000000010";
                        f_reg(362) <= "00100000000111010000000000000000";
                        f_reg(363) <= "00010100111101010000000000111100";
                        f_reg(364) <= "10101111101001110000011111100000";
                        f_reg(365) <= "10001100000111010000100001000000";
                        f_reg(366) <= "00011111101000000000000000000011";
                        f_reg(367) <= "00100000000111010000000000111100";
                        f_reg(368) <= "00010000000000000000000000000010";
                        f_reg(369) <= "00100000000111010000000000000000";
                        f_reg(370) <= "00010101000101100000000000110101";
                        f_reg(371) <= "10101111101010000000011111100100";
                        f_reg(372) <= "10001100000111010000100001000000";
                        f_reg(373) <= "00011111101000000000000000000011";
                        f_reg(374) <= "00100000000111010000000000111100";
                        f_reg(375) <= "00010000000000000000000000000010";
                        f_reg(376) <= "00100000000111010000000000000000";
                        f_reg(377) <= "00010101001101110000000000101110";
                        f_reg(378) <= "10101111101010010000011111101000";
                        f_reg(379) <= "10001100000111010000100001000000";
                        f_reg(380) <= "00011111101000000000000000000011";
                        f_reg(381) <= "00100000000111010000000000111100";
                        f_reg(382) <= "00010000000000000000000000000010";
                        f_reg(383) <= "00100000000111010000000000000000";
                        f_reg(384) <= "00010101010110000000000000100111";
                        f_reg(385) <= "10101111101010100000011111101100";
                        f_reg(386) <= "10001100000111010000100001000000";
                        f_reg(387) <= "00011111101000000000000000000011";
                        f_reg(388) <= "00100000000111010000000000111100";
                        f_reg(389) <= "00010000000000000000000000000010";
                        f_reg(390) <= "00100000000111010000000000000000";
                        f_reg(391) <= "00010101011110010000000000100000";
                        f_reg(392) <= "10101111101010110000011111110000";
                        f_reg(393) <= "10001100000111010000100001000000";
                        f_reg(394) <= "00011111101000000000000000000011";
                        f_reg(395) <= "00100000000111010000000000111100";
                        f_reg(396) <= "00010000000000000000000000000010";
                        f_reg(397) <= "00100000000111010000000000000000";
                        f_reg(398) <= "00010101100110100000000000011001";
                        f_reg(399) <= "10101111101011000000011111110100";
                        f_reg(400) <= "10001100000111010000100001000000";
                        f_reg(401) <= "00011111101000000000000000000011";
                        f_reg(402) <= "00100000000111010000000000111100";
                        f_reg(403) <= "00010000000000000000000000000010";
                        f_reg(404) <= "00100000000111010000000000000000";
                        f_reg(405) <= "00010101101110110000000000010010";
                        f_reg(406) <= "10101111101011010000011111111000";
                        f_reg(407) <= "10001100000111010000100001000000";
                        f_reg(408) <= "00011111101000000000000000000011";
                        f_reg(409) <= "00100000000111010000000000111100";
                        f_reg(410) <= "00010000000000000000000000000010";
                        f_reg(411) <= "00100000000111010000000000000000";
                        f_reg(412) <= "00010101110111000000000000001011";
                        f_reg(413) <= "10101111101011100000011111111100";
                        f_reg(414) <= "10001100000111010000100001000000";
                        f_reg(415) <= "00011111101000000000000000000011";
                        f_reg(416) <= "00100000000111010000000000111100";
                        f_reg(417) <= "00010000000000000000000000000010";
                        f_reg(418) <= "00100000000111010000000000000000";
                        f_reg(419) <= "00010111110111110000000000000100";
                        f_reg(420) <= "10101111101111100000100000000000";
                        f_reg(421) <= "10101100000111010000100001000000";
                        f_reg(422) <= "00010000000000001111111101111011";
                        f_reg(423) <= "10001100000111010000100001000000";
                        f_reg(424) <= "10001111101000010000011111001000";
                        f_reg(425) <= "10001100000111010000100001000000";
                        f_reg(426) <= "10001111101011110000011111001000";
                        f_reg(427) <= "00010100001011111111111111111100";
                        f_reg(428) <= "10001100000111010000100001000000";
                        f_reg(429) <= "10001111101000100000011111001100";
                        f_reg(430) <= "10001100000111010000100001000000";
                        f_reg(431) <= "10001111101100000000011111001100";
                        f_reg(432) <= "00010100010100001111111111111100";
                        f_reg(433) <= "10001100000111010000100001000000";
                        f_reg(434) <= "10001111101000110000011111010000";
                        f_reg(435) <= "10001100000111010000100001000000";
                        f_reg(436) <= "10001111101100010000011111010000";
                        f_reg(437) <= "00010100011100011111111111111100";
                        f_reg(438) <= "10001100000111010000100001000000";
                        f_reg(439) <= "10001111101001000000011111010100";
                        f_reg(440) <= "10001100000111010000100001000000";
                        f_reg(441) <= "10001111101100100000011111010100";
                        f_reg(442) <= "00010100100100101111111111111100";
                        f_reg(443) <= "10001100000111010000100001000000";
                        f_reg(444) <= "10001111101001010000011111011000";
                        f_reg(445) <= "10001100000111010000100001000000";
                        f_reg(446) <= "10001111101100110000011111011000";
                        f_reg(447) <= "00010100101100111111111111111100";
                        f_reg(448) <= "10001100000111010000100001000000";
                        f_reg(449) <= "10001111101001100000011111011100";
                        f_reg(450) <= "10001100000111010000100001000000";
                        f_reg(451) <= "10001111101101000000011111011100";
                        f_reg(452) <= "00010100110101001111111111111100";
                        f_reg(453) <= "10001100000111010000100001000000";
                        f_reg(454) <= "10001111101001110000011111100000";
                        f_reg(455) <= "10001100000111010000100001000000";
                        f_reg(456) <= "10001111101101010000011111100000";
                        f_reg(457) <= "00010100111101011111111111111100";
                        f_reg(458) <= "10001100000111010000100001000000";
                        f_reg(459) <= "10001111101010000000011111100100";
                        f_reg(460) <= "10001100000111010000100001000000";
                        f_reg(461) <= "10001111101101100000011111100100";
                        f_reg(462) <= "00010101000101101111111111111100";
                        f_reg(463) <= "10001100000111010000100001000000";
                        f_reg(464) <= "10001111101010010000011111101000";
                        f_reg(465) <= "10001100000111010000100001000000";
                        f_reg(466) <= "10001111101101110000011111101000";
                        f_reg(467) <= "00010101001101111111111111111100";
                        f_reg(468) <= "10001100000111010000100001000000";
                        f_reg(469) <= "10001111101010100000011111101100";
                        f_reg(470) <= "10001100000111010000100001000000";
                        f_reg(471) <= "10001111101110000000011111101100";
                        f_reg(472) <= "00010101010110001111111111111100";
                        f_reg(473) <= "10001100000111010000100001000000";
                        f_reg(474) <= "10001111101010110000011111110000";
                        f_reg(475) <= "10001100000111010000100001000000";
                        f_reg(476) <= "10001111101110010000011111110000";
                        f_reg(477) <= "00010101011110011111111111111100";
                        f_reg(478) <= "10001100000111010000100001000000";
                        f_reg(479) <= "10001111101011000000011111110100";
                        f_reg(480) <= "10001100000111010000100001000000";
                        f_reg(481) <= "10001111101110100000011111110100";
                        f_reg(482) <= "00010101100110101111111111111100";
                        f_reg(483) <= "10001100000111010000100001000000";
                        f_reg(484) <= "10001111101011010000011111111000";
                        f_reg(485) <= "10001100000111010000100001000000";
                        f_reg(486) <= "10001111101110110000011111111000";
                        f_reg(487) <= "00010101101110111111111111111100";
                        f_reg(488) <= "10001100000111010000100001000000";
                        f_reg(489) <= "10001111101011100000011111111100";
                        f_reg(490) <= "10001100000111010000100001000000";
                        f_reg(491) <= "10001111101111000000011111111100";
                        f_reg(492) <= "00010101110111001111111111111100";
                        f_reg(493) <= "10001100000111010000100001000000";
                        f_reg(494) <= "10001111101111100000100000000000";
                        f_reg(495) <= "10001100000111010000100001000000";
                        f_reg(496) <= "10001111101111110000100000000000";
                        f_reg(497) <= "00010111110111111111111111111100";
                        f_reg(498) <= "00010000000000001111111100101111";
                        f_reg(499) <= "00000000000000000000000000000000";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000001111100111";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                        f_reg(534) <= "00000000000000000000000000000000";
                        f_reg(535) <= "00000000000000000000000000000000";
                        f_reg(536) <= "00000000000000000000000000000000";
                        f_reg(537) <= "00000000000000000000000000000000";
                        f_reg(538) <= "00000000000000000000000000000000";
                        f_reg(539) <= "00000000000000000000000000000000";
                        f_reg(540) <= "00000000000000000000000000000000";
                        f_reg(541) <= "00000000000000000000000000000000";
                        f_reg(542) <= "00000000000000000000000000000000";
                        f_reg(543) <= "00000000000000000000000000000000";
                        f_reg(544) <= "00000000000000000000000000000000";
                        f_reg(545) <= "00000000000000000000000000000000";
                        f_reg(546) <= "00000000000000000000000000000000";
                        f_reg(547) <= "00000000000000000000000000000000";
                        f_reg(548) <= "00000000000000000000000000000000";
                        f_reg(549) <= "00000000000000000000000000000000";
                        f_reg(550) <= "00000000000000000000000000000000";
                        f_reg(551) <= "00000000000000000000000000000000";
                        f_reg(552) <= "00000000000000000000000000000000";
                        f_reg(553) <= "00000000000000000000000000000000";
                        f_reg(554) <= "00000000000000000000000000000000";
                        f_reg(555) <= "00000000000000000000000000000000";
                        f_reg(556) <= "00000000000000000000000000000000";
                        f_reg(557) <= "00000000000000000000000000000000";
                        f_reg(558) <= "00000000000000000000000000000000";
                        f_reg(559) <= "00000000000000000000000000000000";
                        f_reg(560) <= "00000000000000000000000000000000";
                        f_reg(561) <= "00000000000000000000000000000000";
                        f_reg(562) <= "00000000000000000000000000000000";
                        f_reg(563) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test49_Reg_COMBINED;
