--| Test79_Reg_COMBINED.vhd
--| Author: Nicolas Hamilton using write_TMR_VHDL_MEMULATOR.m
--| Created:  18 April 2019 at 15:13:37
--| Emulate the behaviour of a 32-bit addressable memory.  Uses incoming
--| address to determine which instruction to return next.  For write
--| operations, a single internal register will retain the value of i_data
--| until it is overwritten by the next write operation.  Write operations
--| occur when i_write_enable is '1'.
--|
--| INPUTS:
--| i_clk            - clock input
--| i_reset          - reset input
--| i_address	    - address
--| i_read_enable    - enable read
--| i_write_enable   - enable write
--| i_data           - input data
--| i_ack            - acknowlegement that error buffer has received an error
--|
--| OUTPUTS:
--| o_data           - output data
--| o_MEM_READY      - signal is 1 when read/write operation is complete
--| o_DONE           - signal is 1 when the instruction set is completed
--| o_DONE2          - Copy of o_DONE that is sent to a different output pin
--| o_error_detected - signal is 1 when an error has been detected
--| o_error          - indicates the type and location of the error
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test79_Reg_COMBINED is
   port (i_clk             : in  std_logic;
         i_reset           : in  std_logic;
         i_address         : in  std_logic_vector(31 downto 0);
         i_read_enable     : in  std_logic;
         i_write_enable    : in  std_logic;
         i_data            : in  std_logic_vector(31 downto 0);
         i_ack             : in  std_logic;
         o_data            : out std_logic_vector(31 downto 0);
         o_MEM_READY       : out std_logic;
         o_DONE            : out std_logic;
         o_DONE2           : out std_logic;
         o_error_detected  : out std_logic;
         o_error           : out std_logic_vector(39 downto 0));
end Test79_Reg_COMBINED;

architecture a_Test79_Reg_COMBINED of Test79_Reg_COMBINED is
   --| Declare types to store memory addresses and values to store
   type addresses is array (1 to 534) of std_logic_vector (32-1 downto 0);
   type registers is array (1 to 534) of std_logic_vector (32-1 downto 0);

   --| Declare Signals
   -- Registers to delay the ready signal and ensure address is ready to be sampled by the processor
   signal f_MEM_READY : std_logic := '0';
   signal ff_MEM_READY : std_logic := '0';

   -- Registers to store the last value of i_read and i_write
   signal f_read : std_logic := '0';
   signal f_write : std_logic := '0';

   -- Register for data output
   signal f_data : std_logic_vector(31 downto 0) := (others => '0');

   -- Register for the o_DONE output
   signal f_done : std_logic := '0';

   -- Registers for program counter and program flow errors
   signal f_sw_instr       : std_logic := '0'; -- Store word instruction Flag
   signal f_lw_instr       : std_logic := '0'; -- Load word instruction Flag
   signal f_br_instr       : std_logic := '0'; -- Banch instruction flag
   signal f_last_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of last instruction
   signal f_next_address   : std_logic_vector(31 downto 0) := (others => '0'); -- Address of next instruction
   signal f_sw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to store word on write
   signal f_lw_address     : std_logic_vector(31 downto 0) := (others => '0'); -- Address to load word on read
   signal f_branch_address : std_logic_vector(31 downto 0) := (others => '0'); -- Address to branch to on branch instruction

   -- Registers for recovery error detection
   signal f_timeout_flag : std_logic := '0';
   signal f_recovery_flag : std_logic := '0';

   -- Register for timeout error detection
   signal f_clk_count : unsigned(9 downto 0) := (others => '0');

   -- Registers for error outputs
   signal f_error_detected : std_logic := '0'; -- Signal error detection to error buffer
   signal f_error_flag     : std_logic := '0'; -- If error detected while another is being acknowledged by the error buffer
   signal f_error          : std_logic_vector(39 downto 0) := (others => '0'); -- Error data to send to error buffer

   -- Initialize constant for timeout error detection
   constant k_timeout1 : unsigned(9 downto 0) := "0000010100";
   constant k_timeout2 : unsigned(9 downto 0) := "1111101000";

   -- Initialize constants for error types
   constant k_errA : std_logic_vector(7 downto 0) := "01000001";
   constant k_errB : std_logic_vector(7 downto 0) := "01000010";
   constant k_errC : std_logic_vector(7 downto 0) := "01000011";
   constant k_errD : std_logic_vector(7 downto 0) := "01000100";
   constant k_errE : std_logic_vector(7 downto 0) := "01000101";
   constant k_errF : std_logic_vector(7 downto 0) := "01000110";
   constant k_errG : std_logic_vector(7 downto 0) := "01000111";
   constant k_errH : std_logic_vector(7 downto 0) := "01001000";
   constant k_errI : std_logic_vector(7 downto 0) := "01001001";
   constant k_errJ : std_logic_vector(7 downto 0) := "01001010";
   constant k_errK : std_logic_vector(7 downto 0) := "01001011";
   constant k_errX : std_logic_vector(7 downto 0) := "01011000";

   -- Initialize constants for instruction opcodes
   constant k_sw_opcode : std_logic_vector (5 downto 0) := "101011";
   constant k_lw_opcode : std_logic_vector (5 downto 0) := "100011";
   constant k_bgez_bltz_opcode : std_logic_vector (5 downto 0) := "000001";
   constant k_beq_opcode : std_logic_vector (5 downto 0) := "000100";
   constant k_bne_opcode : std_logic_vector (5 downto 0) := "000101";
   constant k_blez_opcode : std_logic_vector (5 downto 0) := "000110";
   constant k_bgtz_opcode : std_logic_vector (5 downto 0) := "000111";

   -- Initialize additional constants
   constant k_zero2 : std_logic_vector (1 downto 0) := (others => '0');
   constant k_zero14 : std_logic_vector (13 downto 0) := (others => '0');
   constant k_zero16 : std_logic_vector (15 downto 0) := (others => '0');
   constant k_ones14 : std_logic_vector (13 downto 0) := (others => '1');
   constant k_four32 : std_logic_vector (31 downto 0) := "00000000000000000000000000000100";

   -- Initialize addresses
   constant k_prog : addresses := (-- Instruction Number - Memory Address
      "00000000000000000000000000000000", --    0 -    0
      "00000000000000000000000000000100", --    1 -    4
      "00000000000000000000000000001000", --    2 -    8
      "00000000000000000000000000001100", --    3 -   12
      "00000000000000000000000000010000", --    4 -   16
      "00000000000000000000000000010100", --    5 -   20
      "00000000000000000000000000011000", --    6 -   24
      "00000000000000000000000000011100", --    7 -   28
      "00000000000000000000000000100000", --    8 -   32
      "00000000000000000000000000100100", --    9 -   36
      "00000000000000000000000000101000", --   10 -   40
      "00000000000000000000000000101100", --   11 -   44
      "00000000000000000000000000110000", --   12 -   48
      "00000000000000000000000000110100", --   13 -   52
      "00000000000000000000000000111000", --   14 -   56
      "00000000000000000000000000111100", --   15 -   60
      "00000000000000000000000001000000", --   16 -   64
      "00000000000000000000000001000100", --   17 -   68
      "00000000000000000000000001001000", --   18 -   72
      "00000000000000000000000001001100", --   19 -   76
      "00000000000000000000000001010000", --   20 -   80
      "00000000000000000000000001010100", --   21 -   84
      "00000000000000000000000001011000", --   22 -   88
      "00000000000000000000000001011100", --   23 -   92
      "00000000000000000000000001100000", --   24 -   96
      "00000000000000000000000001100100", --   25 -  100
      "00000000000000000000000001101000", --   26 -  104
      "00000000000000000000000001101100", --   27 -  108
      "00000000000000000000000001110000", --   28 -  112
      "00000000000000000000000001110100", --   29 -  116
      "00000000000000000000000001111000", --   30 -  120
      "00000000000000000000000001111100", --   31 -  124
      "00000000000000000000000010000000", --   32 -  128
      "00000000000000000000000010000100", --   33 -  132
      "00000000000000000000000010001000", --   34 -  136
      "00000000000000000000000010001100", --   35 -  140
      "00000000000000000000000010010000", --   36 -  144
      "00000000000000000000000010010100", --   37 -  148
      "00000000000000000000000010011000", --   38 -  152
      "00000000000000000000000010011100", --   39 -  156
      "00000000000000000000000010100000", --   40 -  160
      "00000000000000000000000010100100", --   41 -  164
      "00000000000000000000000010101000", --   42 -  168
      "00000000000000000000000010101100", --   43 -  172
      "00000000000000000000000010110000", --   44 -  176
      "00000000000000000000000010110100", --   45 -  180
      "00000000000000000000000010111000", --   46 -  184
      "00000000000000000000000010111100", --   47 -  188
      "00000000000000000000000011000000", --   48 -  192
      "00000000000000000000000011000100", --   49 -  196
      "00000000000000000000000011001000", --   50 -  200
      "00000000000000000000000011001100", --   51 -  204
      "00000000000000000000000011010000", --   52 -  208
      "00000000000000000000000011010100", --   53 -  212
      "00000000000000000000000011011000", --   54 -  216
      "00000000000000000000000011011100", --   55 -  220
      "00000000000000000000000011100000", --   56 -  224
      "00000000000000000000000011100100", --   57 -  228
      "00000000000000000000000011101000", --   58 -  232
      "00000000000000000000000011101100", --   59 -  236
      "00000000000000000000000011110000", --   60 -  240
      "00000000000000000000000011110100", --   61 -  244
      "00000000000000000000000011111000", --   62 -  248
      "00000000000000000000000011111100", --   63 -  252
      "00000000000000000000000100000000", --   64 -  256
      "00000000000000000000000100000100", --   65 -  260
      "00000000000000000000000100001000", --   66 -  264
      "00000000000000000000000100001100", --   67 -  268
      "00000000000000000000000100010000", --   68 -  272
      "00000000000000000000000100010100", --   69 -  276
      "00000000000000000000000100011000", --   70 -  280
      "00000000000000000000000100011100", --   71 -  284
      "00000000000000000000000100100000", --   72 -  288
      "00000000000000000000000100100100", --   73 -  292
      "00000000000000000000000100101000", --   74 -  296
      "00000000000000000000000100101100", --   75 -  300
      "00000000000000000000000100110000", --   76 -  304
      "00000000000000000000000100110100", --   77 -  308
      "00000000000000000000000100111000", --   78 -  312
      "00000000000000000000000100111100", --   79 -  316
      "00000000000000000000000101000000", --   80 -  320
      "00000000000000000000000101000100", --   81 -  324
      "00000000000000000000000101001000", --   82 -  328
      "00000000000000000000000101001100", --   83 -  332
      "00000000000000000000000101010000", --   84 -  336
      "00000000000000000000000101010100", --   85 -  340
      "00000000000000000000000101011000", --   86 -  344
      "00000000000000000000000101011100", --   87 -  348
      "00000000000000000000000101100000", --   88 -  352
      "00000000000000000000000101100100", --   89 -  356
      "00000000000000000000000101101000", --   90 -  360
      "00000000000000000000000101101100", --   91 -  364
      "00000000000000000000000101110000", --   92 -  368
      "00000000000000000000000101110100", --   93 -  372
      "00000000000000000000000101111000", --   94 -  376
      "00000000000000000000000101111100", --   95 -  380
      "00000000000000000000000110000000", --   96 -  384
      "00000000000000000000000110000100", --   97 -  388
      "00000000000000000000000110001000", --   98 -  392
      "00000000000000000000000110001100", --   99 -  396
      "00000000000000000000000110010000", --  100 -  400
      "00000000000000000000000110010100", --  101 -  404
      "00000000000000000000000110011000", --  102 -  408
      "00000000000000000000000110011100", --  103 -  412
      "00000000000000000000000110100000", --  104 -  416
      "00000000000000000000000110100100", --  105 -  420
      "00000000000000000000000110101000", --  106 -  424
      "00000000000000000000000110101100", --  107 -  428
      "00000000000000000000000110110000", --  108 -  432
      "00000000000000000000000110110100", --  109 -  436
      "00000000000000000000000110111000", --  110 -  440
      "00000000000000000000000110111100", --  111 -  444
      "00000000000000000000000111000000", --  112 -  448
      "00000000000000000000000111000100", --  113 -  452
      "00000000000000000000000111001000", --  114 -  456
      "00000000000000000000000111001100", --  115 -  460
      "00000000000000000000000111010000", --  116 -  464
      "00000000000000000000000111010100", --  117 -  468
      "00000000000000000000000111011000", --  118 -  472
      "00000000000000000000000111011100", --  119 -  476
      "00000000000000000000000111100000", --  120 -  480
      "00000000000000000000000111100100", --  121 -  484
      "00000000000000000000000111101000", --  122 -  488
      "00000000000000000000000111101100", --  123 -  492
      "00000000000000000000000111110000", --  124 -  496
      "00000000000000000000000111110100", --  125 -  500
      "00000000000000000000000111111000", --  126 -  504
      "00000000000000000000000111111100", --  127 -  508
      "00000000000000000000001000000000", --  128 -  512
      "00000000000000000000001000000100", --  129 -  516
      "00000000000000000000001000001000", --  130 -  520
      "00000000000000000000001000001100", --  131 -  524
      "00000000000000000000001000010000", --  132 -  528
      "00000000000000000000001000010100", --  133 -  532
      "00000000000000000000001000011000", --  134 -  536
      "00000000000000000000001000011100", --  135 -  540
      "00000000000000000000001000100000", --  136 -  544
      "00000000000000000000001000100100", --  137 -  548
      "00000000000000000000001000101000", --  138 -  552
      "00000000000000000000001000101100", --  139 -  556
      "00000000000000000000001000110000", --  140 -  560
      "00000000000000000000001000110100", --  141 -  564
      "00000000000000000000001000111000", --  142 -  568
      "00000000000000000000001000111100", --  143 -  572
      "00000000000000000000001001000000", --  144 -  576
      "00000000000000000000001001000100", --  145 -  580
      "00000000000000000000001001001000", --  146 -  584
      "00000000000000000000001001001100", --  147 -  588
      "00000000000000000000001001010000", --  148 -  592
      "00000000000000000000001001010100", --  149 -  596
      "00000000000000000000001001011000", --  150 -  600
      "00000000000000000000001001011100", --  151 -  604
      "00000000000000000000001001100000", --  152 -  608
      "00000000000000000000001001100100", --  153 -  612
      "00000000000000000000001001101000", --  154 -  616
      "00000000000000000000001001101100", --  155 -  620
      "00000000000000000000001001110000", --  156 -  624
      "00000000000000000000001001110100", --  157 -  628
      "00000000000000000000001001111000", --  158 -  632
      "00000000000000000000001001111100", --  159 -  636
      "00000000000000000000001010000000", --  160 -  640
      "00000000000000000000001010000100", --  161 -  644
      "00000000000000000000001010001000", --  162 -  648
      "00000000000000000000001010001100", --  163 -  652
      "00000000000000000000001010010000", --  164 -  656
      "00000000000000000000001010010100", --  165 -  660
      "00000000000000000000001010011000", --  166 -  664
      "00000000000000000000001010011100", --  167 -  668
      "00000000000000000000001010100000", --  168 -  672
      "00000000000000000000001010100100", --  169 -  676
      "00000000000000000000001010101000", --  170 -  680
      "00000000000000000000001010101100", --  171 -  684
      "00000000000000000000001010110000", --  172 -  688
      "00000000000000000000001010110100", --  173 -  692
      "00000000000000000000001010111000", --  174 -  696
      "00000000000000000000001010111100", --  175 -  700
      "00000000000000000000001011000000", --  176 -  704
      "00000000000000000000001011000100", --  177 -  708
      "00000000000000000000001011001000", --  178 -  712
      "00000000000000000000001011001100", --  179 -  716
      "00000000000000000000001011010000", --  180 -  720
      "00000000000000000000001011010100", --  181 -  724
      "00000000000000000000001011011000", --  182 -  728
      "00000000000000000000001011011100", --  183 -  732
      "00000000000000000000001011100000", --  184 -  736
      "00000000000000000000001011100100", --  185 -  740
      "00000000000000000000001011101000", --  186 -  744
      "00000000000000000000001011101100", --  187 -  748
      "00000000000000000000001011110000", --  188 -  752
      "00000000000000000000001011110100", --  189 -  756
      "00000000000000000000001011111000", --  190 -  760
      "00000000000000000000001011111100", --  191 -  764
      "00000000000000000000001100000000", --  192 -  768
      "00000000000000000000001100000100", --  193 -  772
      "00000000000000000000001100001000", --  194 -  776
      "00000000000000000000001100001100", --  195 -  780
      "00000000000000000000001100010000", --  196 -  784
      "00000000000000000000001100010100", --  197 -  788
      "00000000000000000000001100011000", --  198 -  792
      "00000000000000000000001100011100", --  199 -  796
      "00000000000000000000001100100000", --  200 -  800
      "00000000000000000000001100100100", --  201 -  804
      "00000000000000000000001100101000", --  202 -  808
      "00000000000000000000001100101100", --  203 -  812
      "00000000000000000000001100110000", --  204 -  816
      "00000000000000000000001100110100", --  205 -  820
      "00000000000000000000001100111000", --  206 -  824
      "00000000000000000000001100111100", --  207 -  828
      "00000000000000000000001101000000", --  208 -  832
      "00000000000000000000001101000100", --  209 -  836
      "00000000000000000000001101001000", --  210 -  840
      "00000000000000000000001101001100", --  211 -  844
      "00000000000000000000001101010000", --  212 -  848
      "00000000000000000000001101010100", --  213 -  852
      "00000000000000000000001101011000", --  214 -  856
      "00000000000000000000001101011100", --  215 -  860
      "00000000000000000000001101100000", --  216 -  864
      "00000000000000000000001101100100", --  217 -  868
      "00000000000000000000001101101000", --  218 -  872
      "00000000000000000000001101101100", --  219 -  876
      "00000000000000000000001101110000", --  220 -  880
      "00000000000000000000001101110100", --  221 -  884
      "00000000000000000000001101111000", --  222 -  888
      "00000000000000000000001101111100", --  223 -  892
      "00000000000000000000001110000000", --  224 -  896
      "00000000000000000000001110000100", --  225 -  900
      "00000000000000000000001110001000", --  226 -  904
      "00000000000000000000001110001100", --  227 -  908
      "00000000000000000000001110010000", --  228 -  912
      "00000000000000000000001110010100", --  229 -  916
      "00000000000000000000001110011000", --  230 -  920
      "00000000000000000000001110011100", --  231 -  924
      "00000000000000000000001110100000", --  232 -  928
      "00000000000000000000001110100100", --  233 -  932
      "00000000000000000000001110101000", --  234 -  936
      "00000000000000000000001110101100", --  235 -  940
      "00000000000000000000001110110000", --  236 -  944
      "00000000000000000000001110110100", --  237 -  948
      "00000000000000000000001110111000", --  238 -  952
      "00000000000000000000001110111100", --  239 -  956
      "00000000000000000000001111000000", --  240 -  960
      "00000000000000000000001111000100", --  241 -  964
      "00000000000000000000001111001000", --  242 -  968
      "00000000000000000000001111001100", --  243 -  972
      "00000000000000000000001111010000", --  244 -  976
      "00000000000000000000001111010100", --  245 -  980
      "00000000000000000000001111011000", --  246 -  984
      "00000000000000000000001111011100", --  247 -  988
      "00000000000000000000001111100000", --  248 -  992
      "00000000000000000000001111100100", --  249 -  996
      "00000000000000000000001111101000", --  250 - 1000
      "00000000000000000000001111101100", --  251 - 1004
      "00000000000000000000001111110000", --  252 - 1008
      "00000000000000000000001111110100", --  253 - 1012
      "00000000000000000000001111111000", --  254 - 1016
      "00000000000000000000001111111100", --  255 - 1020
      "00000000000000000000010000000000", --  256 - 1024
      "00000000000000000000010000000100", --  257 - 1028
      "00000000000000000000010000001000", --  258 - 1032
      "00000000000000000000010000001100", --  259 - 1036
      "00000000000000000000010000010000", --  260 - 1040
      "00000000000000000000010000010100", --  261 - 1044
      "00000000000000000000010000011000", --  262 - 1048
      "00000000000000000000010000011100", --  263 - 1052
      "00000000000000000000010000100000", --  264 - 1056
      "00000000000000000000010000100100", --  265 - 1060
      "00000000000000000000010000101000", --  266 - 1064
      "00000000000000000000010000101100", --  267 - 1068
      "00000000000000000000010000110000", --  268 - 1072
      "00000000000000000000010000110100", --  269 - 1076
      "00000000000000000000010000111000", --  270 - 1080
      "00000000000000000000010000111100", --  271 - 1084
      "00000000000000000000010001000000", --  272 - 1088
      "00000000000000000000010001000100", --  273 - 1092
      "00000000000000000000010001001000", --  274 - 1096
      "00000000000000000000010001001100", --  275 - 1100
      "00000000000000000000010001010000", --  276 - 1104
      "00000000000000000000010001010100", --  277 - 1108
      "00000000000000000000010001011000", --  278 - 1112
      "00000000000000000000010001011100", --  279 - 1116
      "00000000000000000000010001100000", --  280 - 1120
      "00000000000000000000010001100100", --  281 - 1124
      "00000000000000000000010001101000", --  282 - 1128
      "00000000000000000000010001101100", --  283 - 1132
      "00000000000000000000010001110000", --  284 - 1136
      "00000000000000000000010001110100", --  285 - 1140
      "00000000000000000000010001111000", --  286 - 1144
      "00000000000000000000010001111100", --  287 - 1148
      "00000000000000000000010010000000", --  288 - 1152
      "00000000000000000000010010000100", --  289 - 1156
      "00000000000000000000010010001000", --  290 - 1160
      "00000000000000000000010010001100", --  291 - 1164
      "00000000000000000000010010010000", --  292 - 1168
      "00000000000000000000010010010100", --  293 - 1172
      "00000000000000000000010010011000", --  294 - 1176
      "00000000000000000000010010011100", --  295 - 1180
      "00000000000000000000010010100000", --  296 - 1184
      "00000000000000000000010010100100", --  297 - 1188
      "00000000000000000000010010101000", --  298 - 1192
      "00000000000000000000010010101100", --  299 - 1196
      "00000000000000000000010010110000", --  300 - 1200
      "00000000000000000000010010110100", --  301 - 1204
      "00000000000000000000010010111000", --  302 - 1208
      "00000000000000000000010010111100", --  303 - 1212
      "00000000000000000000010011000000", --  304 - 1216
      "00000000000000000000010011000100", --  305 - 1220
      "00000000000000000000010011001000", --  306 - 1224
      "00000000000000000000010011001100", --  307 - 1228
      "00000000000000000000010011010000", --  308 - 1232
      "00000000000000000000010011010100", --  309 - 1236
      "00000000000000000000010011011000", --  310 - 1240
      "00000000000000000000010011011100", --  311 - 1244
      "00000000000000000000010011100000", --  312 - 1248
      "00000000000000000000010011100100", --  313 - 1252
      "00000000000000000000010011101000", --  314 - 1256
      "00000000000000000000010011101100", --  315 - 1260
      "00000000000000000000010011110000", --  316 - 1264
      "00000000000000000000010011110100", --  317 - 1268
      "00000000000000000000010011111000", --  318 - 1272
      "00000000000000000000010011111100", --  319 - 1276
      "00000000000000000000010100000000", --  320 - 1280
      "00000000000000000000010100000100", --  321 - 1284
      "00000000000000000000010100001000", --  322 - 1288
      "00000000000000000000010100001100", --  323 - 1292
      "00000000000000000000010100010000", --  324 - 1296
      "00000000000000000000010100010100", --  325 - 1300
      "00000000000000000000010100011000", --  326 - 1304
      "00000000000000000000010100011100", --  327 - 1308
      "00000000000000000000010100100000", --  328 - 1312
      "00000000000000000000010100100100", --  329 - 1316
      "00000000000000000000010100101000", --  330 - 1320
      "00000000000000000000010100101100", --  331 - 1324
      "00000000000000000000010100110000", --  332 - 1328
      "00000000000000000000010100110100", --  333 - 1332
      "00000000000000000000010100111000", --  334 - 1336
      "00000000000000000000010100111100", --  335 - 1340
      "00000000000000000000010101000000", --  336 - 1344
      "00000000000000000000010101000100", --  337 - 1348
      "00000000000000000000010101001000", --  338 - 1352
      "00000000000000000000010101001100", --  339 - 1356
      "00000000000000000000010101010000", --  340 - 1360
      "00000000000000000000010101010100", --  341 - 1364
      "00000000000000000000010101011000", --  342 - 1368
      "00000000000000000000010101011100", --  343 - 1372
      "00000000000000000000010101100000", --  344 - 1376
      "00000000000000000000010101100100", --  345 - 1380
      "00000000000000000000010101101000", --  346 - 1384
      "00000000000000000000010101101100", --  347 - 1388
      "00000000000000000000010101110000", --  348 - 1392
      "00000000000000000000010101110100", --  349 - 1396
      "00000000000000000000010101111000", --  350 - 1400
      "00000000000000000000010101111100", --  351 - 1404
      "00000000000000000000010110000000", --  352 - 1408
      "00000000000000000000010110000100", --  353 - 1412
      "00000000000000000000010110001000", --  354 - 1416
      "00000000000000000000010110001100", --  355 - 1420
      "00000000000000000000010110010000", --  356 - 1424
      "00000000000000000000010110010100", --  357 - 1428
      "00000000000000000000010110011000", --  358 - 1432
      "00000000000000000000010110011100", --  359 - 1436
      "00000000000000000000010110100000", --  360 - 1440
      "00000000000000000000010110100100", --  361 - 1444
      "00000000000000000000010110101000", --  362 - 1448
      "00000000000000000000010110101100", --  363 - 1452
      "00000000000000000000010110110000", --  364 - 1456
      "00000000000000000000010110110100", --  365 - 1460
      "00000000000000000000010110111000", --  366 - 1464
      "00000000000000000000010110111100", --  367 - 1468
      "00000000000000000000010111000000", --  368 - 1472
      "00000000000000000000010111000100", --  369 - 1476
      "00000000000000000000010111001000", --  370 - 1480
      "00000000000000000000010111001100", --  371 - 1484
      "00000000000000000000010111010000", --  372 - 1488
      "00000000000000000000010111010100", --  373 - 1492
      "00000000000000000000010111011000", --  374 - 1496
      "00000000000000000000010111011100", --  375 - 1500
      "00000000000000000000010111100000", --  376 - 1504
      "00000000000000000000010111100100", --  377 - 1508
      "00000000000000000000010111101000", --  378 - 1512
      "00000000000000000000010111101100", --  379 - 1516
      "00000000000000000000010111110000", --  380 - 1520
      "00000000000000000000010111110100", --  381 - 1524
      "00000000000000000000010111111000", --  382 - 1528
      "00000000000000000000010111111100", --  383 - 1532
      "00000000000000000000011000000000", --  384 - 1536
      "00000000000000000000011000000100", --  385 - 1540
      "00000000000000000000011000001000", --  386 - 1544
      "00000000000000000000011000001100", --  387 - 1548
      "00000000000000000000011000010000", --  388 - 1552
      "00000000000000000000011000010100", --  389 - 1556
      "00000000000000000000011000011000", --  390 - 1560
      "00000000000000000000011000011100", --  391 - 1564
      "00000000000000000000011000100000", --  392 - 1568
      "00000000000000000000011000100100", --  393 - 1572
      "00000000000000000000011000101000", --  394 - 1576
      "00000000000000000000011000101100", --  395 - 1580
      "00000000000000000000011000110000", --  396 - 1584
      "00000000000000000000011000110100", --  397 - 1588
      "00000000000000000000011000111000", --  398 - 1592
      "00000000000000000000011000111100", --  399 - 1596
      "00000000000000000000011001000000", --  400 - 1600
      "00000000000000000000011001000100", --  401 - 1604
      "00000000000000000000011001001000", --  402 - 1608
      "00000000000000000000011001001100", --  403 - 1612
      "00000000000000000000011001010000", --  404 - 1616
      "00000000000000000000011001010100", --  405 - 1620
      "00000000000000000000011001011000", --  406 - 1624
      "00000000000000000000011001011100", --  407 - 1628
      "00000000000000000000011001100000", --  408 - 1632
      "00000000000000000000011001100100", --  409 - 1636
      "00000000000000000000011001101000", --  410 - 1640
      "00000000000000000000011001101100", --  411 - 1644
      "00000000000000000000011001110000", --  412 - 1648
      "00000000000000000000011001110100", --  413 - 1652
      "00000000000000000000011001111000", --  414 - 1656
      "00000000000000000000011001111100", --  415 - 1660
      "00000000000000000000011010000000", --  416 - 1664
      "00000000000000000000011010000100", --  417 - 1668
      "00000000000000000000011010001000", --  418 - 1672
      "00000000000000000000011010001100", --  419 - 1676
      "00000000000000000000011010010000", --  420 - 1680
      "00000000000000000000011010010100", --  421 - 1684
      "00000000000000000000011010011000", --  422 - 1688
      "00000000000000000000011010011100", --  423 - 1692
      "00000000000000000000011010100000", --  424 - 1696
      "00000000000000000000011010100100", --  425 - 1700
      "00000000000000000000011010101000", --  426 - 1704
      "00000000000000000000011010101100", --  427 - 1708
      "00000000000000000000011010110000", --  428 - 1712
      "00000000000000000000011010110100", --  429 - 1716
      "00000000000000000000011010111000", --  430 - 1720
      "00000000000000000000011010111100", --  431 - 1724
      "00000000000000000000011011000000", --  432 - 1728
      "00000000000000000000011011000100", --  433 - 1732
      "00000000000000000000011011001000", --  434 - 1736
      "00000000000000000000011011001100", --  435 - 1740
      "00000000000000000000011011010000", --  436 - 1744
      "00000000000000000000011011010100", --  437 - 1748
      "00000000000000000000011011011000", --  438 - 1752
      "00000000000000000000011011011100", --  439 - 1756
      "00000000000000000000011011100000", --  440 - 1760
      "00000000000000000000011011100100", --  441 - 1764
      "00000000000000000000011011101000", --  442 - 1768
      "00000000000000000000011011101100", --  443 - 1772
      "00000000000000000000011011110000", --  444 - 1776
      "00000000000000000000011011110100", --  445 - 1780
      "00000000000000000000011011111000", --  446 - 1784
      "00000000000000000000011011111100", --  447 - 1788
      "00000000000000000000011100000000", --  448 - 1792
      "00000000000000000000011100000100", --  449 - 1796
      "00000000000000000000011100001000", --  450 - 1800
      "00000000000000000000011100001100", --  451 - 1804
      "00000000000000000000011100010000", --  452 - 1808
      "00000000000000000000011100010100", --  453 - 1812
      "00000000000000000000011100011000", --  454 - 1816
      "00000000000000000000011100011100", --  455 - 1820
      "00000000000000000000011100100000", --  456 - 1824
      "00000000000000000000011100100100", --  457 - 1828
      "00000000000000000000011100101000", --  458 - 1832
      "00000000000000000000011100101100", --  459 - 1836
      "00000000000000000000011100110000", --  460 - 1840
      "00000000000000000000011100110100", --  461 - 1844
      "00000000000000000000011100111000", --  462 - 1848
      "00000000000000000000011100111100", --  463 - 1852
      "00000000000000000000011101000000", --  464 - 1856
      "00000000000000000000011101000100", --  465 - 1860
      "00000000000000000000011101001000", --  466 - 1864
      "00000000000000000000011101001100", --  467 - 1868
      "00000000000000000000011101010000", --  468 - 1872
      "00000000000000000000011101010100", --  469 - 1876
      "00000000000000000000011101011000", --  470 - 1880
      "00000000000000000000011101011100", --  471 - 1884
      "00000000000000000000011101100000", --  472 - 1888
      "00000000000000000000011101100100", --  473 - 1892
      "00000000000000000000011101101000", --  474 - 1896
      "00000000000000000000011101101100", --  475 - 1900
      "00000000000000000000011101110000", --  476 - 1904
      "00000000000000000000011101110100", --  477 - 1908
      "00000000000000000000011101111000", --  478 - 1912
      "00000000000000000000011101111100", --  479 - 1916
      "00000000000000000000011110000000", --  480 - 1920
      "00000000000000000000011110000100", --  481 - 1924
      "00000000000000000000011110001000", --  482 - 1928
      "00000000000000000000011110001100", --  483 - 1932
      "00000000000000000000011110010000", --  484 - 1936
      "00000000000000000000011110010100", --  485 - 1940
      "00000000000000000000011110011000", --  486 - 1944
      "00000000000000000000011110011100", --  487 - 1948
      "00000000000000000000011110100000", --  488 - 1952
      "00000000000000000000011110100100", --  489 - 1956
      "00000000000000000000011110101000", --  490 - 1960
      "00000000000000000000011110101100", --  491 - 1964
      "00000000000000000000011110110000", --  492 - 1968
      "00000000000000000000011110110100", --  493 - 1972
      "00000000000000000000011110111000", --  494 - 1976
      "00000000000000000000011110111100", --  495 - 1980
      "00000000000000000000011111000000", --  496 - 1984
      "00000000000000000000011111000100", --  497 - 1988
      "00000000000000000000011111001000", --  498 - 1992
      "00000000000000000000011111001100", --  499 - 1996
      "00000000000000000000011111010000", --  500 - 2000
      "00000000000000000000011111010100", --  501 - 2004
      "00000000000000000000011111011000", --  502 - 2008
      "00000000000000000000011111011100", --  503 - 2012
      "00000000000000000000011111100000", --  504 - 2016
      "00000000000000000000011111100100", --  505 - 2020
      "00000000000000000000011111101000", --  506 - 2024
      "00000000000000000000011111101100", --  507 - 2028
      "00000000000000000000011111110000", --  508 - 2032
      "00000000000000000000011111110100", --  509 - 2036
      "00000000000000000000011111111000", --  510 - 2040
      "00000000000000000000011111111100", --  511 - 2044
      "00000000000000000000100000000000", --  512 - 2048
      "00000000000000000000100000000100", --  513 - 2052
      "00000000000000000000100000001000", --  514 - 2056
      "00000000000000000000100000001100", --  515 - 2060
      "00000000000000000000100000010000", --  516 - 2064
      "00000000000000000000100000010100", --  517 - 2068
      "00000000000000000000100000011000", --  518 - 2072
      "00000000000000000000100000011100", --  519 - 2076
      "00000000000000000000100000100000", --  520 - 2080
      "00000000000000000000100000100100", --  521 - 2084
      "00000000000000000000100000101000", --  522 - 2088
      "00000000000000000000100000101100", --  523 - 2092
      "00000000000000000000100000110000", --  524 - 2096
      "00000000000000000000100000110100", --  525 - 2100
      "00000000000000000000100000111000", --  526 - 2104
      "00000000000000000000100000111100", --  527 - 2108
      "00000000000000000000100001000000", --  528 - 2112
      "00000000000000000000100001000100", --  529 - 2116
      "00000000000000000000100001001000", --  530 - 2120
      "00000000000000000000100001001100", --  531 - 2124
      "00000000000000000000100001010000", --  532 - 2128
      "00000000000000000000100001010100");--  533 - 2132

   --| Initialize values stored in memory
   signal f_reg: registers := (-- Instruction Number - Memory Address
      "00111100000111110000001111100111", --    0 -    0
      "00000000000111111111110000000010", --    1 -    4
      "00111100000000011011010000101011", --    2 -    8
      "00000000001000000001000000101011", --    3 -   12
      "00111000010000111100011011001011", --    4 -   16
      "00000000011000100010000000000100", --    5 -   20
      "00000000001000110010100000101010", --    6 -   24
      "00101100100001100111001010011100", --    7 -   28
      "00101100110001111101001000000111", --    8 -   32
      "00000000111001110100000000100110", --    9 -   36
      "00110100101010010110110010111101", --   10 -   40
      "00000000010001010101000000000110", --   11 -   44
      "00000000000001110101110010000000", --   12 -   48
      "10101100000000110000010000111000", --   13 -   52
      "00000000010010010110000000100010", --   14 -   56
      "00000000100000000110100000100101", --   15 -   60
      "00110100000011100111011010100001", --   16 -   64
      "00000001100011010111100000101010", --   17 -   68
      "00000001000011111000000000000110", --   18 -   72
      "00000000010011111000100000100110", --   19 -   76
      "00111100000100100010010111000101", --   20 -   80
      "00000000000001011001110101000000", --   21 -   84
      "00000001101011101010000000101011", --   22 -   88
      "00000000010000101010100000100011", --   23 -   92
      "00000000011011100111000000000100", --   24 -   96
      "00100100011101101001011111000111", --   25 -  100
      "00000010110100001011100000000110", --   26 -  104
      "00110010100110000111111001111001", --   27 -  108
      "00000000100110001100100000100011", --   28 -  112
      "10101100000100100000010000111100", --   29 -  116
      "00000001001101011101000000000111", --   30 -  120
      "00100111010110111101000101111101", --   31 -  124
      "00000011000010101110000000100101", --   32 -  128
      "00110100101111010110100111001000", --   33 -  132
      "10101100000111000000010001000000", --   34 -  136
      "00000010111001101111000000000110", --   35 -  140
      "00000011010101100000100000100101", --   36 -  144
      "10101100000111000000010001000100", --   37 -  148
      "00110011110011001010100010100010", --   38 -  152
      "00000001001111010100000000101010", --   39 -  156
      "00000001100001000010000000100110", --   40 -  160
      "00000001110110110111100000101010", --   41 -  164
      "00000001011100010001000000100011", --   42 -  168
      "00000000000011000001100101000010", --   43 -  172
      "00000001000100111000000000100010", --   44 -  176
      "00000000100001111010000000100110", --   45 -  180
      "00000000010011011001000000100001", --   46 -  184
      "00000000111000011010100000000100", --   47 -  188
      "00101100011010100110000110110111", --   48 -  192
      "00000010101110010010100000100111", --   49 -  196
      "00000000000000000000000000000000", --   50 -  200
      "00101110011001100101110000011101", --   51 -  204
      "00000010010001011011100000000100", --   52 -  208
      "00101011011110100111010011110100", --   53 -  212
      "00000000000011111011001110000010", --   54 -  216
      "00000000000000000000000000000000", --   55 -  220
      "10101100000100110000010001001000", --   56 -  224
      "00110011010111001111100100000000", --   57 -  228
      "00000010111101000100100000100111", --   58 -  232
      "00111100000111011011111101100111", --   59 -  236
      "00000001010100000111000000000111", --   60 -  240
      "00000001110001100101100000100100", --   61 -  244
      "00000000000000000000000000000000", --   62 -  248
      "10101100000010110000010001001100", --   63 -  252
      "00000010110101101000100000100110", --   64 -  256
      "10101100000111100000010001010000", --   65 -  260
      "00000000000000000110011000000000", --   66 -  264
      "00100111101010000010000000101001", --   67 -  268
      "00000010001110000010000000100111", --   68 -  272
      "00000001101010000001000000000110", --   69 -  276
      "00000000000000000000000000000000", --   70 -  280
      "00000001100111000000100000100110", --   71 -  284
      "00000000010000010011100000000100", --   72 -  288
      "00000000000000000000000000000000", --   73 -  292
      "10101100000010010000010001010100", --   74 -  296
      "10101100000001110000010001011000", --   75 -  300
      "10101100000001000000010001011100", --   76 -  304
      "00100011111111111111111111111111", --   77 -  308
      "00011111111000001111111110110100", --   78 -  312
      "00010000000000000000000111000110", --   79 -  316
      "00111100000111100000001111100111", --   80 -  320
      "00111100000111110000001111100111", --   81 -  324
      "00000000000111101111010000000010", --   82 -  328
      "00000000000111111111110000000010", --   83 -  332
      "00111100000000011011010000101011", --   84 -  336
      "00111100000011111011010000101011", --   85 -  340
      "00000000001000000001000000101011", --   86 -  344
      "00000001111000001000000000101011", --   87 -  348
      "00111000010000111100011011001011", --   88 -  352
      "00111010000100011100011011001011", --   89 -  356
      "00000000011000100010000000000100", --   90 -  360
      "00000010001100001001000000000100", --   91 -  364
      "00000000001000110010100000101010", --   92 -  368
      "00000001111100011001100000101010", --   93 -  372
      "00101100100001100111001010011100", --   94 -  376
      "00101110010101000111001010011100", --   95 -  380
      "00101100110001111101001000000111", --   96 -  384
      "00101110100101011101001000000111", --   97 -  388
      "00000000111001110100000000100110", --   98 -  392
      "00000010101101011011000000100110", --   99 -  396
      "00110100101010010110110010111101", --  100 -  400
      "00110110011101110110110010111101", --  101 -  404
      "00000000010001010101000000000110", --  102 -  408
      "00000010000100111100000000000110", --  103 -  412
      "00000000000001110101110010000000", --  104 -  416
      "00000000000101011100110010000000", --  105 -  420
      "00010100011100010000000100011110", --  106 -  424
      "10101100000000110000010000111000", --  107 -  428
      "00000000010010010110000000100010", --  108 -  432
      "00000010000101111101000000100010", --  109 -  436
      "00000000100000000110100000100101", --  110 -  440
      "00000010010000001101100000100101", --  111 -  444
      "00110100000011100111011010100001", --  112 -  448
      "00110100000111000111011010100001", --  113 -  452
      "00000001100011010000100000101010", --  114 -  456
      "00000011010110110111100000101010", --  115 -  460
      "00000001000000010110000000000110", --  116 -  464
      "00000010110011111101000000000110", --  117 -  468
      "00000000010000010100000000100110", --  118 -  472
      "00000010000011111011000000100110", --  119 -  476
      "00111100000000010010010111000101", --  120 -  480
      "00111100000011110010010111000101", --  121 -  484
      "00010101101110110000000100001110", --  122 -  488
      "10101100000011010000010001100000", --  123 -  492
      "00000000000001010110110101000000", --  124 -  496
      "00000000000100111101110101000000", --  125 -  500
      "00010101101110110000000100001010", --  126 -  504
      "10101100000011010000010001100100", --  127 -  508
      "10001100000011010000010001100000", --  128 -  512
      "10001100000110110000010001100000", --  129 -  516
      "00010101101110111111111111111110", --  130 -  520
      "00010100111101010000000100000101", --  131 -  524
      "10101100000001110000010001101000", --  132 -  528
      "00000001101011100011100000101011", --  133 -  532
      "00000011011111001010100000101011", --  134 -  536
      "00010101101110110000000100000001", --  135 -  540
      "10101100000011010000010001101100", --  136 -  544
      "00000000010000100110100000100011", --  137 -  548
      "00000010000100001101100000100011", --  138 -  552
      "00000000011011100111000000000100", --  139 -  556
      "00000010001111001110000000000100", --  140 -  560
      "00100100011000101001011111000111", --  141 -  564
      "00100110001100001001011111000111", --  142 -  568
      "00000000010011000001100000000110", --  143 -  572
      "00000010000110101000100000000110", --  144 -  576
      "00110000111011000111111001111001", --  145 -  580
      "00110010101110100111111001111001", --  146 -  584
      "00000000100011000011100000100011", --  147 -  588
      "00000010010110101010100000100011", --  148 -  592
      "00010100001011110000000011110011", --  149 -  596
      "10101100000000010000010000111100", --  150 -  600
      "00000001001011010000100000000111", --  151 -  604
      "00000010111110110111100000000111", --  152 -  608
      "00100100001011011101000101111101", --  153 -  612
      "00100101111110111101000101111101", --  154 -  616
      "00010101101110110000000011101101", --  155 -  620
      "10101100000011010000010001110000", --  156 -  624
      "00000001100010100110100000100101", --  157 -  628
      "00000011010110001101100000100101", --  158 -  632
      "00110100101010100110100111001000", --  159 -  636
      "00110110011110000110100111001000", --  160 -  640
      "00010101101110110000000011100111", --  161 -  644
      "10101100000011010000010001000000", --  162 -  648
      "00000000011001100010100000000110", --  163 -  652
      "00000010001101001001100000000110", --  164 -  656
      "00000000001000100011000000100101", --  165 -  660
      "00000001111100001010000000100101", --  166 -  664
      "00010101101110110000000011100001", --  167 -  668
      "10101100000011010000010001000100", --  168 -  672
      "00110000101000111010100010100010", --  169 -  676
      "00110010011100011010100010100010", --  170 -  680
      "00000001001010100000100000101010", --  171 -  684
      "00000010111110000111100000101010", --  172 -  688
      "00000000011001000010000000100110", --  173 -  692
      "00000010001100101001000000100110", --  174 -  696
      "10001100000000100000010001110000", --  175 -  700
      "10001100000100000000010001110000", --  176 -  704
      "00010100010100001111111111111110", --  177 -  708
      "00000001110000100110100000101010", --  178 -  712
      "00000011100100001101100000101010", --  179 -  716
      "00000001011010000100100000100011", --  180 -  720
      "00000011001101101011100000100011", --  181 -  724
      "00000000000000110101000101000010", --  182 -  728
      "00000000000100011100000101000010", --  183 -  732
      "10001100000011100000010001100100", --  184 -  736
      "10001100000111000000010001100100", --  185 -  740
      "00010101110111001111111111111110", --  186 -  744
      "00000000001011100101100000100010", --  187 -  748
      "00000001111111001100100000100010", --  188 -  752
      "10001100000010000000010001101000", --  189 -  756
      "10001100000101100000010001101000", --  190 -  760
      "00010101000101101111111111111110", --  191 -  764
      "00000000100010000001100000100110", --  192 -  768
      "00000010010101101000100000100110", --  193 -  772
      "10001100000000010000010001101100", --  194 -  776
      "10001100000011110000010001101100", --  195 -  780
      "00010100001011111111111111111110", --  196 -  784
      "00000001001000010010000000100001", --  197 -  788
      "00000010111011111001000000100001", --  198 -  792
      "00000001000001100100100000000100", --  199 -  796
      "00000010110101001011100000000100", --  200 -  800
      "00101101010001100110000110110111", --  201 -  804
      "00101111000101000110000110110111", --  202 -  808
      "00000001001001110100000000100111", --  203 -  812
      "00000010111101011011000000100111", --  204 -  816
      "00000000000000000000000000000000", --  205 -  820
      "00000000000000000000000000000000", --  206 -  824
      "00101101110010100101110000011101", --  207 -  828
      "00101111100110000101110000011101", --  208 -  832
      "00000000100010000100100000000100", --  209 -  836
      "00000010010101101011100000000100", --  210 -  840
      "00101000010001110111010011110100", --  211 -  844
      "00101010000101010111010011110100", --  212 -  848
      "00000000000011010100001110000010", --  213 -  852
      "00000000000110111011001110000010", --  214 -  856
      "00000000000000000000000000000000", --  215 -  860
      "00000000000000000000000000000000", --  216 -  864
      "00010101110111000000000010101111", --  217 -  868
      "10101100000011100000010001001000", --  218 -  872
      "00110000111001001111100100000000", --  219 -  876
      "00110010101100101111100100000000", --  220 -  880
      "00000001001000110001000000100111", --  221 -  884
      "00000010111100011000000000100111", --  222 -  888
      "00111100000011011011111101100111", --  223 -  892
      "00111100000110111011111101100111", --  224 -  896
      "00000000110010110111000000000111", --  225 -  900
      "00000010100110011110000000000111", --  226 -  904
      "00000001110010100011100000100100", --  227 -  908
      "00000011100110001010100000100100", --  228 -  912
      "00000000000000000000000000000000", --  229 -  916
      "00000000000000000000000000000000", --  230 -  920
      "00010100111101010000000010100001", --  231 -  924
      "10101100000001110000010001001100", --  232 -  928
      "00000001000010000100100000100110", --  233 -  932
      "00000010110101101011100000100110", --  234 -  936
      "00010100101100110000000010011101", --  235 -  940
      "10101100000001010000010001010000", --  236 -  944
      "00000000000000000001111000000000", --  237 -  948
      "00000000000000001000111000000000", --  238 -  952
      "00100101101010110010000000101001", --  239 -  956
      "00100111011110010010000000101001", --  240 -  960
      "00000001001011000011000000100111", --  241 -  964
      "00000010111110101010000000100111", --  242 -  968
      "00000000001010110111000000000110", --  243 -  972
      "00000001111110011110000000000110", --  244 -  976
      "00000000000000000000000000000000", --  245 -  980
      "00000000000000000000000000000000", --  246 -  984
      "00000000011001000101000000100110", --  247 -  988
      "00000010001100101100000000100110", --  248 -  992
      "00000001110010100011100000000100", --  249 -  996
      "00000011100110001010100000000100", --  250 - 1000
      "00000000000000000000000000000000", --  251 - 1004
      "00000000000000000000000000000000", --  252 - 1008
      "00010100010100000000000010001011", --  253 - 1012
      "10101100000000100000010001010100", --  254 - 1016
      "00010100111101010000000010001001", --  255 - 1020
      "10101100000001110000010001011000", --  256 - 1024
      "00010100110101000000000010000111", --  257 - 1028
      "10101100000001100000010001011100", --  258 - 1032
      "00100011110111011111111100000110", --  259 - 1036
      "00010011101000000000000000011001", --  260 - 1040
      "00100011110111011111111000001100", --  261 - 1044
      "00010011101000000000000000010111", --  262 - 1048
      "00100011110111011111110100010010", --  263 - 1052
      "00010011101000000000000000010101", --  264 - 1056
      "00100011110111101111111111111111", --  265 - 1060
      "00100011111111111111111111111111", --  266 - 1064
      "00010111110111110000000001111101", --  267 - 1068
      "00011111111000001111111101001000", --  268 - 1072
      "00010000000000000000000100001000", --  269 - 1076
      "00000000000000000000000000000000", --  270 - 1080
      "00000000000000000000000000000000", --  271 - 1084
      "00000000000000000000000000000000", --  272 - 1088
      "00000000000000000000000000000000", --  273 - 1092
      "00000000000000000000000000000000", --  274 - 1096
      "00000000000000000000000000000000", --  275 - 1100
      "00000000000000000000000000000000", --  276 - 1104
      "00000000000000000000000000000000", --  277 - 1108
      "00000000000000000000000000000000", --  278 - 1112
      "00000000000000000000000000000000", --  279 - 1116
      "00000000000000000000000000000000", --  280 - 1120
      "00000000000000000000000000000000", --  281 - 1124
      "00000000000000000000000000000000", --  282 - 1128
      "00000000000000000000000000000000", --  283 - 1132
      "00000000000000000000000000000000", --  284 - 1136
      "10001100000111010000011111001000", --  285 - 1140
      "00011111101000000000000000000011", --  286 - 1144
      "00100000000111010000000000111100", --  287 - 1148
      "00010000000000000000000000000010", --  288 - 1152
      "00100000000111010000000000000000", --  289 - 1156
      "00010100001011110000000001100110", --  290 - 1160
      "10101111101000010000011101010000", --  291 - 1164
      "10001100000111010000011111001000", --  292 - 1168
      "00011111101000000000000000000011", --  293 - 1172
      "00100000000111010000000000111100", --  294 - 1176
      "00010000000000000000000000000010", --  295 - 1180
      "00100000000111010000000000000000", --  296 - 1184
      "00010100010100000000000001011111", --  297 - 1188
      "10101111101000100000011101010100", --  298 - 1192
      "10001100000111010000011111001000", --  299 - 1196
      "00011111101000000000000000000011", --  300 - 1200
      "00100000000111010000000000111100", --  301 - 1204
      "00010000000000000000000000000010", --  302 - 1208
      "00100000000111010000000000000000", --  303 - 1212
      "00010100011100010000000001011000", --  304 - 1216
      "10101111101000110000011101011000", --  305 - 1220
      "10001100000111010000011111001000", --  306 - 1224
      "00011111101000000000000000000011", --  307 - 1228
      "00100000000111010000000000111100", --  308 - 1232
      "00010000000000000000000000000010", --  309 - 1236
      "00100000000111010000000000000000", --  310 - 1240
      "00010100100100100000000001010001", --  311 - 1244
      "10101111101001000000011101011100", --  312 - 1248
      "10001100000111010000011111001000", --  313 - 1252
      "00011111101000000000000000000011", --  314 - 1256
      "00100000000111010000000000111100", --  315 - 1260
      "00010000000000000000000000000010", --  316 - 1264
      "00100000000111010000000000000000", --  317 - 1268
      "00010100101100110000000001001010", --  318 - 1272
      "10101111101001010000011101100000", --  319 - 1276
      "10001100000111010000011111001000", --  320 - 1280
      "00011111101000000000000000000011", --  321 - 1284
      "00100000000111010000000000111100", --  322 - 1288
      "00010000000000000000000000000010", --  323 - 1292
      "00100000000111010000000000000000", --  324 - 1296
      "00010100110101000000000001000011", --  325 - 1300
      "10101111101001100000011101100100", --  326 - 1304
      "10001100000111010000011111001000", --  327 - 1308
      "00011111101000000000000000000011", --  328 - 1312
      "00100000000111010000000000111100", --  329 - 1316
      "00010000000000000000000000000010", --  330 - 1320
      "00100000000111010000000000000000", --  331 - 1324
      "00010100111101010000000000111100", --  332 - 1328
      "10101111101001110000011101101000", --  333 - 1332
      "10001100000111010000011111001000", --  334 - 1336
      "00011111101000000000000000000011", --  335 - 1340
      "00100000000111010000000000111100", --  336 - 1344
      "00010000000000000000000000000010", --  337 - 1348
      "00100000000111010000000000000000", --  338 - 1352
      "00010101000101100000000000110101", --  339 - 1356
      "10101111101010000000011101101100", --  340 - 1360
      "10001100000111010000011111001000", --  341 - 1364
      "00011111101000000000000000000011", --  342 - 1368
      "00100000000111010000000000111100", --  343 - 1372
      "00010000000000000000000000000010", --  344 - 1376
      "00100000000111010000000000000000", --  345 - 1380
      "00010101001101110000000000101110", --  346 - 1384
      "10101111101010010000011101110000", --  347 - 1388
      "10001100000111010000011111001000", --  348 - 1392
      "00011111101000000000000000000011", --  349 - 1396
      "00100000000111010000000000111100", --  350 - 1400
      "00010000000000000000000000000010", --  351 - 1404
      "00100000000111010000000000000000", --  352 - 1408
      "00010101010110000000000000100111", --  353 - 1412
      "10101111101010100000011101110100", --  354 - 1416
      "10001100000111010000011111001000", --  355 - 1420
      "00011111101000000000000000000011", --  356 - 1424
      "00100000000111010000000000111100", --  357 - 1428
      "00010000000000000000000000000010", --  358 - 1432
      "00100000000111010000000000000000", --  359 - 1436
      "00010101011110010000000000100000", --  360 - 1440
      "10101111101010110000011101111000", --  361 - 1444
      "10001100000111010000011111001000", --  362 - 1448
      "00011111101000000000000000000011", --  363 - 1452
      "00100000000111010000000000111100", --  364 - 1456
      "00010000000000000000000000000010", --  365 - 1460
      "00100000000111010000000000000000", --  366 - 1464
      "00010101100110100000000000011001", --  367 - 1468
      "10101111101011000000011101111100", --  368 - 1472
      "10001100000111010000011111001000", --  369 - 1476
      "00011111101000000000000000000011", --  370 - 1480
      "00100000000111010000000000111100", --  371 - 1484
      "00010000000000000000000000000010", --  372 - 1488
      "00100000000111010000000000000000", --  373 - 1492
      "00010101101110110000000000010010", --  374 - 1496
      "10101111101011010000011110000000", --  375 - 1500
      "10001100000111010000011111001000", --  376 - 1504
      "00011111101000000000000000000011", --  377 - 1508
      "00100000000111010000000000111100", --  378 - 1512
      "00010000000000000000000000000010", --  379 - 1516
      "00100000000111010000000000000000", --  380 - 1520
      "00010101110111000000000000001011", --  381 - 1524
      "10101111101011100000011110000100", --  382 - 1528
      "10001100000111010000011111001000", --  383 - 1532
      "00011111101000000000000000000011", --  384 - 1536
      "00100000000111010000000000111100", --  385 - 1540
      "00010000000000000000000000000010", --  386 - 1544
      "00100000000111010000000000000000", --  387 - 1548
      "00010111110111110000000000000100", --  388 - 1552
      "10101111101111100000011110001000", --  389 - 1556
      "10101100000111010000011111001000", --  390 - 1560
      "00010000000000001111111110000010", --  391 - 1564
      "10001100000111010000011111001000", --  392 - 1568
      "10001111101000010000011101010000", --  393 - 1572
      "10001100000111010000011111001000", --  394 - 1576
      "10001111101011110000011101010000", --  395 - 1580
      "00010100001011111111111111111100", --  396 - 1584
      "10001100000111010000011111001000", --  397 - 1588
      "10001111101000100000011101010100", --  398 - 1592
      "10001100000111010000011111001000", --  399 - 1596
      "10001111101100000000011101010100", --  400 - 1600
      "00010100010100001111111111111100", --  401 - 1604
      "10001100000111010000011111001000", --  402 - 1608
      "10001111101000110000011101011000", --  403 - 1612
      "10001100000111010000011111001000", --  404 - 1616
      "10001111101100010000011101011000", --  405 - 1620
      "00010100011100011111111111111100", --  406 - 1624
      "10001100000111010000011111001000", --  407 - 1628
      "10001111101001000000011101011100", --  408 - 1632
      "10001100000111010000011111001000", --  409 - 1636
      "10001111101100100000011101011100", --  410 - 1640
      "00010100100100101111111111111100", --  411 - 1644
      "10001100000111010000011111001000", --  412 - 1648
      "10001111101001010000011101100000", --  413 - 1652
      "10001100000111010000011111001000", --  414 - 1656
      "10001111101100110000011101100000", --  415 - 1660
      "00010100101100111111111111111100", --  416 - 1664
      "10001100000111010000011111001000", --  417 - 1668
      "10001111101001100000011101100100", --  418 - 1672
      "10001100000111010000011111001000", --  419 - 1676
      "10001111101101000000011101100100", --  420 - 1680
      "00010100110101001111111111111100", --  421 - 1684
      "10001100000111010000011111001000", --  422 - 1688
      "10001111101001110000011101101000", --  423 - 1692
      "10001100000111010000011111001000", --  424 - 1696
      "10001111101101010000011101101000", --  425 - 1700
      "00010100111101011111111111111100", --  426 - 1704
      "10001100000111010000011111001000", --  427 - 1708
      "10001111101010000000011101101100", --  428 - 1712
      "10001100000111010000011111001000", --  429 - 1716
      "10001111101101100000011101101100", --  430 - 1720
      "00010101000101101111111111111100", --  431 - 1724
      "10001100000111010000011111001000", --  432 - 1728
      "10001111101010010000011101110000", --  433 - 1732
      "10001100000111010000011111001000", --  434 - 1736
      "10001111101101110000011101110000", --  435 - 1740
      "00010101001101111111111111111100", --  436 - 1744
      "10001100000111010000011111001000", --  437 - 1748
      "10001111101010100000011101110100", --  438 - 1752
      "10001100000111010000011111001000", --  439 - 1756
      "10001111101110000000011101110100", --  440 - 1760
      "00010101010110001111111111111100", --  441 - 1764
      "10001100000111010000011111001000", --  442 - 1768
      "10001111101010110000011101111000", --  443 - 1772
      "10001100000111010000011111001000", --  444 - 1776
      "10001111101110010000011101111000", --  445 - 1780
      "00010101011110011111111111111100", --  446 - 1784
      "10001100000111010000011111001000", --  447 - 1788
      "10001111101011000000011101111100", --  448 - 1792
      "10001100000111010000011111001000", --  449 - 1796
      "10001111101110100000011101111100", --  450 - 1800
      "00010101100110101111111111111100", --  451 - 1804
      "10001100000111010000011111001000", --  452 - 1808
      "10001111101011010000011110000000", --  453 - 1812
      "10001100000111010000011111001000", --  454 - 1816
      "10001111101110110000011110000000", --  455 - 1820
      "00010101101110111111111111111100", --  456 - 1824
      "10001100000111010000011111001000", --  457 - 1828
      "10001111101011100000011110000100", --  458 - 1832
      "10001100000111010000011111001000", --  459 - 1836
      "10001111101111000000011110000100", --  460 - 1840
      "00010101110111001111111111111100", --  461 - 1844
      "10001100000111010000011111001000", --  462 - 1848
      "10001111101111100000011110001000", --  463 - 1852
      "10001100000111010000011111001000", --  464 - 1856
      "10001111101111110000011110001000", --  465 - 1860
      "00010111110111111111111111111100", --  466 - 1864
      "00010000000000001111111100110110", --  467 - 1868
      "00000000000000000000000000000000", --  468 - 1872
      "00000000000000000000000000000000", --  469 - 1876
      "00000000000000000000000000000000", --  470 - 1880
      "00000000000000000000000000000000", --  471 - 1884
      "00000000000000000000000000000000", --  472 - 1888
      "00000000000000000000000000000000", --  473 - 1892
      "00000000000000000000000000000000", --  474 - 1896
      "00000000000000000000000000000000", --  475 - 1900
      "00000000000000000000000000000000", --  476 - 1904
      "00000000000000000000000000000000", --  477 - 1908
      "00000000000000000000000000000000", --  478 - 1912
      "00000000000000000000000000000000", --  479 - 1916
      "00000000000000000000000000000000", --  480 - 1920
      "00000000000000000000000000000000", --  481 - 1924
      "00000000000000000000000000000000", --  482 - 1928
      "00000000000000000000000000000000", --  483 - 1932
      "00000000000000000000000000000000", --  484 - 1936
      "00000000000000000000000000000000", --  485 - 1940
      "00000000000000000000000000000000", --  486 - 1944
      "00000000000000000000000000000000", --  487 - 1948
      "00000000000000000000000000000000", --  488 - 1952
      "00000000000000000000000000000000", --  489 - 1956
      "00000000000000000000000000000000", --  490 - 1960
      "00000000000000000000000000000000", --  491 - 1964
      "00000000000000000000000000000000", --  492 - 1968
      "00000000000000000000000000000000", --  493 - 1972
      "00000000000000000000000000000000", --  494 - 1976
      "00000000000000000000000000000000", --  495 - 1980
      "00000000000000000000000000000000", --  496 - 1984
      "00000000000000000000000000000000", --  497 - 1988
      "00000000000000000000001111100111", --  498 - 1992
      "00000000000000000000000000000000", --  499 - 1996
      "00000000000000000000000000000000", --  500 - 2000
      "00000000000000000000000000000000", --  501 - 2004
      "00000000000000000000000000000000", --  502 - 2008
      "00000000000000000000000000000000", --  503 - 2012
      "00000000000000000000000000000000", --  504 - 2016
      "00000000000000000000000000000000", --  505 - 2020
      "00000000000000000000000000000000", --  506 - 2024
      "00000000000000000000000000000000", --  507 - 2028
      "00000000000000000000000000000000", --  508 - 2032
      "00000000000000000000000000000000", --  509 - 2036
      "00000000000000000000000000000000", --  510 - 2040
      "00000000000000000000000000000000", --  511 - 2044
      "00000000000000000000000000000000", --  512 - 2048
      "00000000000000000000000000000000", --  513 - 2052
      "00000000000000000000000000000000", --  514 - 2056
      "00000000000000000000000000000000", --  515 - 2060
      "00000000000000000000000000000000", --  516 - 2064
      "00000000000000000000000000000000", --  517 - 2068
      "00000000000000000000000000000000", --  518 - 2072
      "00000000000000000000000000000000", --  519 - 2076
      "00000000000000000000000000000000", --  520 - 2080
      "00000000000000000000000000000000", --  521 - 2084
      "00000000000000000000000000000000", --  522 - 2088
      "00000000000000000000000000000000", --  523 - 2092
      "00000000000000000000000000000000", --  524 - 2096
      "00000000000000000000000000000000", --  525 - 2100
      "00000000000000000000000000000000", --  526 - 2104
      "00000000000000000000000000000000", --  527 - 2108
      "00000000000000000000000000000000", --  528 - 2112
      "00000000000000000000000000000000", --  529 - 2116
      "00000000000000000000000000000000", --  530 - 2120
      "00000000000000000000000000000000", --  531 - 2124
      "00000000000000000000000000000000", --  532 - 2128
      "00000000000000000000000000000000");--  533 - 2132

begin
   -- Assign output signals
   o_MEM_READY <= ff_MEM_READY;
   o_DONE <= f_DONE;
   o_DONE2 <= f_DONE;
   o_error <= f_error;
   o_error_detected <= f_error_detected;

   mem_read_process : process (i_clk, i_reset, i_read_enable)
   begin
      o_data <= f_data;
      -- When the reset signal is asserted
      if (i_reset = '1') then
         f_done <= '0';
         f_data <= (others => '0');
         f_MEM_READY <= '0';
         ff_MEM_READY <= '0';
         f_read <= '0';
         f_write <= '0';
         f_sw_instr <= '0';
         f_lw_instr <= '0';
         f_br_instr <= '0';
         f_last_address <= (others => '0');
         f_next_address <= (others => '0');
         f_sw_address <= (others => '0');
         f_lw_address <= (others => '0');
         f_branch_address <= (others => '0');
         f_error_detected <= '0';
         f_error_flag <= '0';
         f_error <= (others => '0');
         f_clk_count <= (others => '0');
         f_timeout_flag <= '0';
         f_recovery_flag <= '0';
         f_reg(1) <= "00111100000111110000001111100111";
         f_reg(2) <= "00000000000111111111110000000010";
         f_reg(3) <= "00111100000000011011010000101011";
         f_reg(4) <= "00000000001000000001000000101011";
         f_reg(5) <= "00111000010000111100011011001011";
         f_reg(6) <= "00000000011000100010000000000100";
         f_reg(7) <= "00000000001000110010100000101010";
         f_reg(8) <= "00101100100001100111001010011100";
         f_reg(9) <= "00101100110001111101001000000111";
         f_reg(10) <= "00000000111001110100000000100110";
         f_reg(11) <= "00110100101010010110110010111101";
         f_reg(12) <= "00000000010001010101000000000110";
         f_reg(13) <= "00000000000001110101110010000000";
         f_reg(14) <= "10101100000000110000010000111000";
         f_reg(15) <= "00000000010010010110000000100010";
         f_reg(16) <= "00000000100000000110100000100101";
         f_reg(17) <= "00110100000011100111011010100001";
         f_reg(18) <= "00000001100011010111100000101010";
         f_reg(19) <= "00000001000011111000000000000110";
         f_reg(20) <= "00000000010011111000100000100110";
         f_reg(21) <= "00111100000100100010010111000101";
         f_reg(22) <= "00000000000001011001110101000000";
         f_reg(23) <= "00000001101011101010000000101011";
         f_reg(24) <= "00000000010000101010100000100011";
         f_reg(25) <= "00000000011011100111000000000100";
         f_reg(26) <= "00100100011101101001011111000111";
         f_reg(27) <= "00000010110100001011100000000110";
         f_reg(28) <= "00110010100110000111111001111001";
         f_reg(29) <= "00000000100110001100100000100011";
         f_reg(30) <= "10101100000100100000010000111100";
         f_reg(31) <= "00000001001101011101000000000111";
         f_reg(32) <= "00100111010110111101000101111101";
         f_reg(33) <= "00000011000010101110000000100101";
         f_reg(34) <= "00110100101111010110100111001000";
         f_reg(35) <= "10101100000111000000010001000000";
         f_reg(36) <= "00000010111001101111000000000110";
         f_reg(37) <= "00000011010101100000100000100101";
         f_reg(38) <= "10101100000111000000010001000100";
         f_reg(39) <= "00110011110011001010100010100010";
         f_reg(40) <= "00000001001111010100000000101010";
         f_reg(41) <= "00000001100001000010000000100110";
         f_reg(42) <= "00000001110110110111100000101010";
         f_reg(43) <= "00000001011100010001000000100011";
         f_reg(44) <= "00000000000011000001100101000010";
         f_reg(45) <= "00000001000100111000000000100010";
         f_reg(46) <= "00000000100001111010000000100110";
         f_reg(47) <= "00000000010011011001000000100001";
         f_reg(48) <= "00000000111000011010100000000100";
         f_reg(49) <= "00101100011010100110000110110111";
         f_reg(50) <= "00000010101110010010100000100111";
         f_reg(51) <= "00000000000000000000000000000000";
         f_reg(52) <= "00101110011001100101110000011101";
         f_reg(53) <= "00000010010001011011100000000100";
         f_reg(54) <= "00101011011110100111010011110100";
         f_reg(55) <= "00000000000011111011001110000010";
         f_reg(56) <= "00000000000000000000000000000000";
         f_reg(57) <= "10101100000100110000010001001000";
         f_reg(58) <= "00110011010111001111100100000000";
         f_reg(59) <= "00000010111101000100100000100111";
         f_reg(60) <= "00111100000111011011111101100111";
         f_reg(61) <= "00000001010100000111000000000111";
         f_reg(62) <= "00000001110001100101100000100100";
         f_reg(63) <= "00000000000000000000000000000000";
         f_reg(64) <= "10101100000010110000010001001100";
         f_reg(65) <= "00000010110101101000100000100110";
         f_reg(66) <= "10101100000111100000010001010000";
         f_reg(67) <= "00000000000000000110011000000000";
         f_reg(68) <= "00100111101010000010000000101001";
         f_reg(69) <= "00000010001110000010000000100111";
         f_reg(70) <= "00000001101010000001000000000110";
         f_reg(71) <= "00000000000000000000000000000000";
         f_reg(72) <= "00000001100111000000100000100110";
         f_reg(73) <= "00000000010000010011100000000100";
         f_reg(74) <= "00000000000000000000000000000000";
         f_reg(75) <= "10101100000010010000010001010100";
         f_reg(76) <= "10101100000001110000010001011000";
         f_reg(77) <= "10101100000001000000010001011100";
         f_reg(78) <= "00100011111111111111111111111111";
         f_reg(79) <= "00011111111000001111111110110100";
         f_reg(80) <= "00010000000000000000000111000110";
         f_reg(81) <= "00111100000111100000001111100111";
         f_reg(82) <= "00111100000111110000001111100111";
         f_reg(83) <= "00000000000111101111010000000010";
         f_reg(84) <= "00000000000111111111110000000010";
         f_reg(85) <= "00111100000000011011010000101011";
         f_reg(86) <= "00111100000011111011010000101011";
         f_reg(87) <= "00000000001000000001000000101011";
         f_reg(88) <= "00000001111000001000000000101011";
         f_reg(89) <= "00111000010000111100011011001011";
         f_reg(90) <= "00111010000100011100011011001011";
         f_reg(91) <= "00000000011000100010000000000100";
         f_reg(92) <= "00000010001100001001000000000100";
         f_reg(93) <= "00000000001000110010100000101010";
         f_reg(94) <= "00000001111100011001100000101010";
         f_reg(95) <= "00101100100001100111001010011100";
         f_reg(96) <= "00101110010101000111001010011100";
         f_reg(97) <= "00101100110001111101001000000111";
         f_reg(98) <= "00101110100101011101001000000111";
         f_reg(99) <= "00000000111001110100000000100110";
         f_reg(100) <= "00000010101101011011000000100110";
         f_reg(101) <= "00110100101010010110110010111101";
         f_reg(102) <= "00110110011101110110110010111101";
         f_reg(103) <= "00000000010001010101000000000110";
         f_reg(104) <= "00000010000100111100000000000110";
         f_reg(105) <= "00000000000001110101110010000000";
         f_reg(106) <= "00000000000101011100110010000000";
         f_reg(107) <= "00010100011100010000000100011110";
         f_reg(108) <= "10101100000000110000010000111000";
         f_reg(109) <= "00000000010010010110000000100010";
         f_reg(110) <= "00000010000101111101000000100010";
         f_reg(111) <= "00000000100000000110100000100101";
         f_reg(112) <= "00000010010000001101100000100101";
         f_reg(113) <= "00110100000011100111011010100001";
         f_reg(114) <= "00110100000111000111011010100001";
         f_reg(115) <= "00000001100011010000100000101010";
         f_reg(116) <= "00000011010110110111100000101010";
         f_reg(117) <= "00000001000000010110000000000110";
         f_reg(118) <= "00000010110011111101000000000110";
         f_reg(119) <= "00000000010000010100000000100110";
         f_reg(120) <= "00000010000011111011000000100110";
         f_reg(121) <= "00111100000000010010010111000101";
         f_reg(122) <= "00111100000011110010010111000101";
         f_reg(123) <= "00010101101110110000000100001110";
         f_reg(124) <= "10101100000011010000010001100000";
         f_reg(125) <= "00000000000001010110110101000000";
         f_reg(126) <= "00000000000100111101110101000000";
         f_reg(127) <= "00010101101110110000000100001010";
         f_reg(128) <= "10101100000011010000010001100100";
         f_reg(129) <= "10001100000011010000010001100000";
         f_reg(130) <= "10001100000110110000010001100000";
         f_reg(131) <= "00010101101110111111111111111110";
         f_reg(132) <= "00010100111101010000000100000101";
         f_reg(133) <= "10101100000001110000010001101000";
         f_reg(134) <= "00000001101011100011100000101011";
         f_reg(135) <= "00000011011111001010100000101011";
         f_reg(136) <= "00010101101110110000000100000001";
         f_reg(137) <= "10101100000011010000010001101100";
         f_reg(138) <= "00000000010000100110100000100011";
         f_reg(139) <= "00000010000100001101100000100011";
         f_reg(140) <= "00000000011011100111000000000100";
         f_reg(141) <= "00000010001111001110000000000100";
         f_reg(142) <= "00100100011000101001011111000111";
         f_reg(143) <= "00100110001100001001011111000111";
         f_reg(144) <= "00000000010011000001100000000110";
         f_reg(145) <= "00000010000110101000100000000110";
         f_reg(146) <= "00110000111011000111111001111001";
         f_reg(147) <= "00110010101110100111111001111001";
         f_reg(148) <= "00000000100011000011100000100011";
         f_reg(149) <= "00000010010110101010100000100011";
         f_reg(150) <= "00010100001011110000000011110011";
         f_reg(151) <= "10101100000000010000010000111100";
         f_reg(152) <= "00000001001011010000100000000111";
         f_reg(153) <= "00000010111110110111100000000111";
         f_reg(154) <= "00100100001011011101000101111101";
         f_reg(155) <= "00100101111110111101000101111101";
         f_reg(156) <= "00010101101110110000000011101101";
         f_reg(157) <= "10101100000011010000010001110000";
         f_reg(158) <= "00000001100010100110100000100101";
         f_reg(159) <= "00000011010110001101100000100101";
         f_reg(160) <= "00110100101010100110100111001000";
         f_reg(161) <= "00110110011110000110100111001000";
         f_reg(162) <= "00010101101110110000000011100111";
         f_reg(163) <= "10101100000011010000010001000000";
         f_reg(164) <= "00000000011001100010100000000110";
         f_reg(165) <= "00000010001101001001100000000110";
         f_reg(166) <= "00000000001000100011000000100101";
         f_reg(167) <= "00000001111100001010000000100101";
         f_reg(168) <= "00010101101110110000000011100001";
         f_reg(169) <= "10101100000011010000010001000100";
         f_reg(170) <= "00110000101000111010100010100010";
         f_reg(171) <= "00110010011100011010100010100010";
         f_reg(172) <= "00000001001010100000100000101010";
         f_reg(173) <= "00000010111110000111100000101010";
         f_reg(174) <= "00000000011001000010000000100110";
         f_reg(175) <= "00000010001100101001000000100110";
         f_reg(176) <= "10001100000000100000010001110000";
         f_reg(177) <= "10001100000100000000010001110000";
         f_reg(178) <= "00010100010100001111111111111110";
         f_reg(179) <= "00000001110000100110100000101010";
         f_reg(180) <= "00000011100100001101100000101010";
         f_reg(181) <= "00000001011010000100100000100011";
         f_reg(182) <= "00000011001101101011100000100011";
         f_reg(183) <= "00000000000000110101000101000010";
         f_reg(184) <= "00000000000100011100000101000010";
         f_reg(185) <= "10001100000011100000010001100100";
         f_reg(186) <= "10001100000111000000010001100100";
         f_reg(187) <= "00010101110111001111111111111110";
         f_reg(188) <= "00000000001011100101100000100010";
         f_reg(189) <= "00000001111111001100100000100010";
         f_reg(190) <= "10001100000010000000010001101000";
         f_reg(191) <= "10001100000101100000010001101000";
         f_reg(192) <= "00010101000101101111111111111110";
         f_reg(193) <= "00000000100010000001100000100110";
         f_reg(194) <= "00000010010101101000100000100110";
         f_reg(195) <= "10001100000000010000010001101100";
         f_reg(196) <= "10001100000011110000010001101100";
         f_reg(197) <= "00010100001011111111111111111110";
         f_reg(198) <= "00000001001000010010000000100001";
         f_reg(199) <= "00000010111011111001000000100001";
         f_reg(200) <= "00000001000001100100100000000100";
         f_reg(201) <= "00000010110101001011100000000100";
         f_reg(202) <= "00101101010001100110000110110111";
         f_reg(203) <= "00101111000101000110000110110111";
         f_reg(204) <= "00000001001001110100000000100111";
         f_reg(205) <= "00000010111101011011000000100111";
         f_reg(206) <= "00000000000000000000000000000000";
         f_reg(207) <= "00000000000000000000000000000000";
         f_reg(208) <= "00101101110010100101110000011101";
         f_reg(209) <= "00101111100110000101110000011101";
         f_reg(210) <= "00000000100010000100100000000100";
         f_reg(211) <= "00000010010101101011100000000100";
         f_reg(212) <= "00101000010001110111010011110100";
         f_reg(213) <= "00101010000101010111010011110100";
         f_reg(214) <= "00000000000011010100001110000010";
         f_reg(215) <= "00000000000110111011001110000010";
         f_reg(216) <= "00000000000000000000000000000000";
         f_reg(217) <= "00000000000000000000000000000000";
         f_reg(218) <= "00010101110111000000000010101111";
         f_reg(219) <= "10101100000011100000010001001000";
         f_reg(220) <= "00110000111001001111100100000000";
         f_reg(221) <= "00110010101100101111100100000000";
         f_reg(222) <= "00000001001000110001000000100111";
         f_reg(223) <= "00000010111100011000000000100111";
         f_reg(224) <= "00111100000011011011111101100111";
         f_reg(225) <= "00111100000110111011111101100111";
         f_reg(226) <= "00000000110010110111000000000111";
         f_reg(227) <= "00000010100110011110000000000111";
         f_reg(228) <= "00000001110010100011100000100100";
         f_reg(229) <= "00000011100110001010100000100100";
         f_reg(230) <= "00000000000000000000000000000000";
         f_reg(231) <= "00000000000000000000000000000000";
         f_reg(232) <= "00010100111101010000000010100001";
         f_reg(233) <= "10101100000001110000010001001100";
         f_reg(234) <= "00000001000010000100100000100110";
         f_reg(235) <= "00000010110101101011100000100110";
         f_reg(236) <= "00010100101100110000000010011101";
         f_reg(237) <= "10101100000001010000010001010000";
         f_reg(238) <= "00000000000000000001111000000000";
         f_reg(239) <= "00000000000000001000111000000000";
         f_reg(240) <= "00100101101010110010000000101001";
         f_reg(241) <= "00100111011110010010000000101001";
         f_reg(242) <= "00000001001011000011000000100111";
         f_reg(243) <= "00000010111110101010000000100111";
         f_reg(244) <= "00000000001010110111000000000110";
         f_reg(245) <= "00000001111110011110000000000110";
         f_reg(246) <= "00000000000000000000000000000000";
         f_reg(247) <= "00000000000000000000000000000000";
         f_reg(248) <= "00000000011001000101000000100110";
         f_reg(249) <= "00000010001100101100000000100110";
         f_reg(250) <= "00000001110010100011100000000100";
         f_reg(251) <= "00000011100110001010100000000100";
         f_reg(252) <= "00000000000000000000000000000000";
         f_reg(253) <= "00000000000000000000000000000000";
         f_reg(254) <= "00010100010100000000000010001011";
         f_reg(255) <= "10101100000000100000010001010100";
         f_reg(256) <= "00010100111101010000000010001001";
         f_reg(257) <= "10101100000001110000010001011000";
         f_reg(258) <= "00010100110101000000000010000111";
         f_reg(259) <= "10101100000001100000010001011100";
         f_reg(260) <= "00100011110111011111111100000110";
         f_reg(261) <= "00010011101000000000000000011001";
         f_reg(262) <= "00100011110111011111111000001100";
         f_reg(263) <= "00010011101000000000000000010111";
         f_reg(264) <= "00100011110111011111110100010010";
         f_reg(265) <= "00010011101000000000000000010101";
         f_reg(266) <= "00100011110111101111111111111111";
         f_reg(267) <= "00100011111111111111111111111111";
         f_reg(268) <= "00010111110111110000000001111101";
         f_reg(269) <= "00011111111000001111111101001000";
         f_reg(270) <= "00010000000000000000000100001000";
         f_reg(271) <= "00000000000000000000000000000000";
         f_reg(272) <= "00000000000000000000000000000000";
         f_reg(273) <= "00000000000000000000000000000000";
         f_reg(274) <= "00000000000000000000000000000000";
         f_reg(275) <= "00000000000000000000000000000000";
         f_reg(276) <= "00000000000000000000000000000000";
         f_reg(277) <= "00000000000000000000000000000000";
         f_reg(278) <= "00000000000000000000000000000000";
         f_reg(279) <= "00000000000000000000000000000000";
         f_reg(280) <= "00000000000000000000000000000000";
         f_reg(281) <= "00000000000000000000000000000000";
         f_reg(282) <= "00000000000000000000000000000000";
         f_reg(283) <= "00000000000000000000000000000000";
         f_reg(284) <= "00000000000000000000000000000000";
         f_reg(285) <= "00000000000000000000000000000000";
         f_reg(286) <= "10001100000111010000011111001000";
         f_reg(287) <= "00011111101000000000000000000011";
         f_reg(288) <= "00100000000111010000000000111100";
         f_reg(289) <= "00010000000000000000000000000010";
         f_reg(290) <= "00100000000111010000000000000000";
         f_reg(291) <= "00010100001011110000000001100110";
         f_reg(292) <= "10101111101000010000011101010000";
         f_reg(293) <= "10001100000111010000011111001000";
         f_reg(294) <= "00011111101000000000000000000011";
         f_reg(295) <= "00100000000111010000000000111100";
         f_reg(296) <= "00010000000000000000000000000010";
         f_reg(297) <= "00100000000111010000000000000000";
         f_reg(298) <= "00010100010100000000000001011111";
         f_reg(299) <= "10101111101000100000011101010100";
         f_reg(300) <= "10001100000111010000011111001000";
         f_reg(301) <= "00011111101000000000000000000011";
         f_reg(302) <= "00100000000111010000000000111100";
         f_reg(303) <= "00010000000000000000000000000010";
         f_reg(304) <= "00100000000111010000000000000000";
         f_reg(305) <= "00010100011100010000000001011000";
         f_reg(306) <= "10101111101000110000011101011000";
         f_reg(307) <= "10001100000111010000011111001000";
         f_reg(308) <= "00011111101000000000000000000011";
         f_reg(309) <= "00100000000111010000000000111100";
         f_reg(310) <= "00010000000000000000000000000010";
         f_reg(311) <= "00100000000111010000000000000000";
         f_reg(312) <= "00010100100100100000000001010001";
         f_reg(313) <= "10101111101001000000011101011100";
         f_reg(314) <= "10001100000111010000011111001000";
         f_reg(315) <= "00011111101000000000000000000011";
         f_reg(316) <= "00100000000111010000000000111100";
         f_reg(317) <= "00010000000000000000000000000010";
         f_reg(318) <= "00100000000111010000000000000000";
         f_reg(319) <= "00010100101100110000000001001010";
         f_reg(320) <= "10101111101001010000011101100000";
         f_reg(321) <= "10001100000111010000011111001000";
         f_reg(322) <= "00011111101000000000000000000011";
         f_reg(323) <= "00100000000111010000000000111100";
         f_reg(324) <= "00010000000000000000000000000010";
         f_reg(325) <= "00100000000111010000000000000000";
         f_reg(326) <= "00010100110101000000000001000011";
         f_reg(327) <= "10101111101001100000011101100100";
         f_reg(328) <= "10001100000111010000011111001000";
         f_reg(329) <= "00011111101000000000000000000011";
         f_reg(330) <= "00100000000111010000000000111100";
         f_reg(331) <= "00010000000000000000000000000010";
         f_reg(332) <= "00100000000111010000000000000000";
         f_reg(333) <= "00010100111101010000000000111100";
         f_reg(334) <= "10101111101001110000011101101000";
         f_reg(335) <= "10001100000111010000011111001000";
         f_reg(336) <= "00011111101000000000000000000011";
         f_reg(337) <= "00100000000111010000000000111100";
         f_reg(338) <= "00010000000000000000000000000010";
         f_reg(339) <= "00100000000111010000000000000000";
         f_reg(340) <= "00010101000101100000000000110101";
         f_reg(341) <= "10101111101010000000011101101100";
         f_reg(342) <= "10001100000111010000011111001000";
         f_reg(343) <= "00011111101000000000000000000011";
         f_reg(344) <= "00100000000111010000000000111100";
         f_reg(345) <= "00010000000000000000000000000010";
         f_reg(346) <= "00100000000111010000000000000000";
         f_reg(347) <= "00010101001101110000000000101110";
         f_reg(348) <= "10101111101010010000011101110000";
         f_reg(349) <= "10001100000111010000011111001000";
         f_reg(350) <= "00011111101000000000000000000011";
         f_reg(351) <= "00100000000111010000000000111100";
         f_reg(352) <= "00010000000000000000000000000010";
         f_reg(353) <= "00100000000111010000000000000000";
         f_reg(354) <= "00010101010110000000000000100111";
         f_reg(355) <= "10101111101010100000011101110100";
         f_reg(356) <= "10001100000111010000011111001000";
         f_reg(357) <= "00011111101000000000000000000011";
         f_reg(358) <= "00100000000111010000000000111100";
         f_reg(359) <= "00010000000000000000000000000010";
         f_reg(360) <= "00100000000111010000000000000000";
         f_reg(361) <= "00010101011110010000000000100000";
         f_reg(362) <= "10101111101010110000011101111000";
         f_reg(363) <= "10001100000111010000011111001000";
         f_reg(364) <= "00011111101000000000000000000011";
         f_reg(365) <= "00100000000111010000000000111100";
         f_reg(366) <= "00010000000000000000000000000010";
         f_reg(367) <= "00100000000111010000000000000000";
         f_reg(368) <= "00010101100110100000000000011001";
         f_reg(369) <= "10101111101011000000011101111100";
         f_reg(370) <= "10001100000111010000011111001000";
         f_reg(371) <= "00011111101000000000000000000011";
         f_reg(372) <= "00100000000111010000000000111100";
         f_reg(373) <= "00010000000000000000000000000010";
         f_reg(374) <= "00100000000111010000000000000000";
         f_reg(375) <= "00010101101110110000000000010010";
         f_reg(376) <= "10101111101011010000011110000000";
         f_reg(377) <= "10001100000111010000011111001000";
         f_reg(378) <= "00011111101000000000000000000011";
         f_reg(379) <= "00100000000111010000000000111100";
         f_reg(380) <= "00010000000000000000000000000010";
         f_reg(381) <= "00100000000111010000000000000000";
         f_reg(382) <= "00010101110111000000000000001011";
         f_reg(383) <= "10101111101011100000011110000100";
         f_reg(384) <= "10001100000111010000011111001000";
         f_reg(385) <= "00011111101000000000000000000011";
         f_reg(386) <= "00100000000111010000000000111100";
         f_reg(387) <= "00010000000000000000000000000010";
         f_reg(388) <= "00100000000111010000000000000000";
         f_reg(389) <= "00010111110111110000000000000100";
         f_reg(390) <= "10101111101111100000011110001000";
         f_reg(391) <= "10101100000111010000011111001000";
         f_reg(392) <= "00010000000000001111111110000010";
         f_reg(393) <= "10001100000111010000011111001000";
         f_reg(394) <= "10001111101000010000011101010000";
         f_reg(395) <= "10001100000111010000011111001000";
         f_reg(396) <= "10001111101011110000011101010000";
         f_reg(397) <= "00010100001011111111111111111100";
         f_reg(398) <= "10001100000111010000011111001000";
         f_reg(399) <= "10001111101000100000011101010100";
         f_reg(400) <= "10001100000111010000011111001000";
         f_reg(401) <= "10001111101100000000011101010100";
         f_reg(402) <= "00010100010100001111111111111100";
         f_reg(403) <= "10001100000111010000011111001000";
         f_reg(404) <= "10001111101000110000011101011000";
         f_reg(405) <= "10001100000111010000011111001000";
         f_reg(406) <= "10001111101100010000011101011000";
         f_reg(407) <= "00010100011100011111111111111100";
         f_reg(408) <= "10001100000111010000011111001000";
         f_reg(409) <= "10001111101001000000011101011100";
         f_reg(410) <= "10001100000111010000011111001000";
         f_reg(411) <= "10001111101100100000011101011100";
         f_reg(412) <= "00010100100100101111111111111100";
         f_reg(413) <= "10001100000111010000011111001000";
         f_reg(414) <= "10001111101001010000011101100000";
         f_reg(415) <= "10001100000111010000011111001000";
         f_reg(416) <= "10001111101100110000011101100000";
         f_reg(417) <= "00010100101100111111111111111100";
         f_reg(418) <= "10001100000111010000011111001000";
         f_reg(419) <= "10001111101001100000011101100100";
         f_reg(420) <= "10001100000111010000011111001000";
         f_reg(421) <= "10001111101101000000011101100100";
         f_reg(422) <= "00010100110101001111111111111100";
         f_reg(423) <= "10001100000111010000011111001000";
         f_reg(424) <= "10001111101001110000011101101000";
         f_reg(425) <= "10001100000111010000011111001000";
         f_reg(426) <= "10001111101101010000011101101000";
         f_reg(427) <= "00010100111101011111111111111100";
         f_reg(428) <= "10001100000111010000011111001000";
         f_reg(429) <= "10001111101010000000011101101100";
         f_reg(430) <= "10001100000111010000011111001000";
         f_reg(431) <= "10001111101101100000011101101100";
         f_reg(432) <= "00010101000101101111111111111100";
         f_reg(433) <= "10001100000111010000011111001000";
         f_reg(434) <= "10001111101010010000011101110000";
         f_reg(435) <= "10001100000111010000011111001000";
         f_reg(436) <= "10001111101101110000011101110000";
         f_reg(437) <= "00010101001101111111111111111100";
         f_reg(438) <= "10001100000111010000011111001000";
         f_reg(439) <= "10001111101010100000011101110100";
         f_reg(440) <= "10001100000111010000011111001000";
         f_reg(441) <= "10001111101110000000011101110100";
         f_reg(442) <= "00010101010110001111111111111100";
         f_reg(443) <= "10001100000111010000011111001000";
         f_reg(444) <= "10001111101010110000011101111000";
         f_reg(445) <= "10001100000111010000011111001000";
         f_reg(446) <= "10001111101110010000011101111000";
         f_reg(447) <= "00010101011110011111111111111100";
         f_reg(448) <= "10001100000111010000011111001000";
         f_reg(449) <= "10001111101011000000011101111100";
         f_reg(450) <= "10001100000111010000011111001000";
         f_reg(451) <= "10001111101110100000011101111100";
         f_reg(452) <= "00010101100110101111111111111100";
         f_reg(453) <= "10001100000111010000011111001000";
         f_reg(454) <= "10001111101011010000011110000000";
         f_reg(455) <= "10001100000111010000011111001000";
         f_reg(456) <= "10001111101110110000011110000000";
         f_reg(457) <= "00010101101110111111111111111100";
         f_reg(458) <= "10001100000111010000011111001000";
         f_reg(459) <= "10001111101011100000011110000100";
         f_reg(460) <= "10001100000111010000011111001000";
         f_reg(461) <= "10001111101111000000011110000100";
         f_reg(462) <= "00010101110111001111111111111100";
         f_reg(463) <= "10001100000111010000011111001000";
         f_reg(464) <= "10001111101111100000011110001000";
         f_reg(465) <= "10001100000111010000011111001000";
         f_reg(466) <= "10001111101111110000011110001000";
         f_reg(467) <= "00010111110111111111111111111100";
         f_reg(468) <= "00010000000000001111111100110110";
         f_reg(469) <= "00000000000000000000000000000000";
         f_reg(470) <= "00000000000000000000000000000000";
         f_reg(471) <= "00000000000000000000000000000000";
         f_reg(472) <= "00000000000000000000000000000000";
         f_reg(473) <= "00000000000000000000000000000000";
         f_reg(474) <= "00000000000000000000000000000000";
         f_reg(475) <= "00000000000000000000000000000000";
         f_reg(476) <= "00000000000000000000000000000000";
         f_reg(477) <= "00000000000000000000000000000000";
         f_reg(478) <= "00000000000000000000000000000000";
         f_reg(479) <= "00000000000000000000000000000000";
         f_reg(480) <= "00000000000000000000000000000000";
         f_reg(481) <= "00000000000000000000000000000000";
         f_reg(482) <= "00000000000000000000000000000000";
         f_reg(483) <= "00000000000000000000000000000000";
         f_reg(484) <= "00000000000000000000000000000000";
         f_reg(485) <= "00000000000000000000000000000000";
         f_reg(486) <= "00000000000000000000000000000000";
         f_reg(487) <= "00000000000000000000000000000000";
         f_reg(488) <= "00000000000000000000000000000000";
         f_reg(489) <= "00000000000000000000000000000000";
         f_reg(490) <= "00000000000000000000000000000000";
         f_reg(491) <= "00000000000000000000000000000000";
         f_reg(492) <= "00000000000000000000000000000000";
         f_reg(493) <= "00000000000000000000000000000000";
         f_reg(494) <= "00000000000000000000000000000000";
         f_reg(495) <= "00000000000000000000000000000000";
         f_reg(496) <= "00000000000000000000000000000000";
         f_reg(497) <= "00000000000000000000000000000000";
         f_reg(498) <= "00000000000000000000000000000000";
         f_reg(499) <= "00000000000000000000001111100111";
         f_reg(500) <= "00000000000000000000000000000000";
         f_reg(501) <= "00000000000000000000000000000000";
         f_reg(502) <= "00000000000000000000000000000000";
         f_reg(503) <= "00000000000000000000000000000000";
         f_reg(504) <= "00000000000000000000000000000000";
         f_reg(505) <= "00000000000000000000000000000000";
         f_reg(506) <= "00000000000000000000000000000000";
         f_reg(507) <= "00000000000000000000000000000000";
         f_reg(508) <= "00000000000000000000000000000000";
         f_reg(509) <= "00000000000000000000000000000000";
         f_reg(510) <= "00000000000000000000000000000000";
         f_reg(511) <= "00000000000000000000000000000000";
         f_reg(512) <= "00000000000000000000000000000000";
         f_reg(513) <= "00000000000000000000000000000000";
         f_reg(514) <= "00000000000000000000000000000000";
         f_reg(515) <= "00000000000000000000000000000000";
         f_reg(516) <= "00000000000000000000000000000000";
         f_reg(517) <= "00000000000000000000000000000000";
         f_reg(518) <= "00000000000000000000000000000000";
         f_reg(519) <= "00000000000000000000000000000000";
         f_reg(520) <= "00000000000000000000000000000000";
         f_reg(521) <= "00000000000000000000000000000000";
         f_reg(522) <= "00000000000000000000000000000000";
         f_reg(523) <= "00000000000000000000000000000000";
         f_reg(524) <= "00000000000000000000000000000000";
         f_reg(525) <= "00000000000000000000000000000000";
         f_reg(526) <= "00000000000000000000000000000000";
         f_reg(527) <= "00000000000000000000000000000000";
         f_reg(528) <= "00000000000000000000000000000000";
         f_reg(529) <= "00000000000000000000000000000000";
         f_reg(530) <= "00000000000000000000000000000000";
         f_reg(531) <= "00000000000000000000000000000000";
         f_reg(532) <= "00000000000000000000000000000000";
         f_reg(533) <= "00000000000000000000000000000000";
      -- At every rising clock edge
      elsif rising_edge(i_clk) then
         if (f_DONE = '0') then
            ff_MEM_READY <= f_MEM_READY;

            -- When attempting to read from memory
            if (i_read_enable = '1') then
               if (f_read = '0') then
                  f_read <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_data <= f_reg(1);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(2);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(3) =>
                        -- LUI R1 -19413
                        f_data <= f_reg(3);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(4) =>
                        -- SLTU R2 R1 R0
                        f_data <= f_reg(4);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(5) =>
                        -- XORI R3 R2 -14645
                        f_data <= f_reg(5);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(6) =>
                        -- SLLV R4 R2 R3
                        f_data <= f_reg(6);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(7) =>
                        -- SLT R5 R1 R3
                        f_data <= f_reg(7);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(8) =>
                        -- SLTIU R6 R4 29340
                        f_data <= f_reg(8);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(9) =>
                        -- SLTIU R7 R6 -11769
                        f_data <= f_reg(9);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(10) =>
                        -- XOR R8 R7 R7
                        f_data <= f_reg(10);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(11) =>
                        -- ORI R9 R5 27837
                        f_data <= f_reg(11);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(12) =>
                        -- SRLV R10 R5 R2
                        f_data <= f_reg(12);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(13) =>
                        -- SLL R11 R7 18
                        f_data <= f_reg(13);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(14) =>
                        -- SW R3 R0 1080
                        f_data <= f_reg(14);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(15) =>
                        -- SUB R12 R2 R9
                        f_data <= f_reg(15);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(16) =>
                        -- OR R13 R4 R0
                        f_data <= f_reg(16);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(17) =>
                        -- ORI R14 R0 30369
                        f_data <= f_reg(17);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(18) =>
                        -- SLT R15 R12 R13
                        f_data <= f_reg(18);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(19) =>
                        -- SRLV R16 R15 R8
                        f_data <= f_reg(19);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(20) =>
                        -- XOR R17 R2 R15
                        f_data <= f_reg(20);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(21) =>
                        -- LUI R18 9669
                        f_data <= f_reg(21);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(22) =>
                        -- SLL R19 R5 21
                        f_data <= f_reg(22);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(23) =>
                        -- SLTU R20 R13 R14
                        f_data <= f_reg(23);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(24) =>
                        -- SUBU R21 R2 R2
                        f_data <= f_reg(24);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(25) =>
                        -- SLLV R14 R14 R3
                        f_data <= f_reg(25);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(26) =>
                        -- ADDIU R22 R3 -26681
                        f_data <= f_reg(26);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(27) =>
                        -- SRLV R23 R16 R22
                        f_data <= f_reg(27);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(28) =>
                        -- ANDI R24 R20 32377
                        f_data <= f_reg(28);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(29) =>
                        -- SUBU R25 R4 R24
                        f_data <= f_reg(29);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(30) =>
                        -- SW R18 R0 1084
                        f_data <= f_reg(30);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(31) =>
                        -- SRAV R26 R21 R9
                        f_data <= f_reg(31);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(32) =>
                        -- ADDIU R27 R26 -11907
                        f_data <= f_reg(32);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(33) =>
                        -- OR R28 R24 R10
                        f_data <= f_reg(33);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(34) =>
                        -- ORI R29 R5 27080
                        f_data <= f_reg(34);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(35) =>
                        -- SW R28 R0 1088
                        f_data <= f_reg(35);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(36) =>
                        -- SRLV R30 R6 R23
                        f_data <= f_reg(36);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(37) =>
                        -- OR R1 R26 R22
                        f_data <= f_reg(37);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(38) =>
                        -- SW R28 R0 1092
                        f_data <= f_reg(38);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(39) =>
                        -- ANDI R12 R30 -22366
                        f_data <= f_reg(39);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(40) =>
                        -- SLT R8 R9 R29
                        f_data <= f_reg(40);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(41) =>
                        -- XOR R4 R12 R4
                        f_data <= f_reg(41);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(42) =>
                        -- SLT R15 R14 R27
                        f_data <= f_reg(42);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(43) =>
                        -- SUBU R2 R11 R17
                        f_data <= f_reg(43);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(44) =>
                        -- SRL R3 R12 5
                        f_data <= f_reg(44);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(45) =>
                        -- SUB R16 R8 R19
                        f_data <= f_reg(45);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(46) =>
                        -- XOR R20 R4 R7
                        f_data <= f_reg(46);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(47) =>
                        -- ADDU R18 R2 R13
                        f_data <= f_reg(47);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(48) =>
                        -- SLLV R21 R1 R7
                        f_data <= f_reg(48);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(49) =>
                        -- SLTIU R10 R3 25015
                        f_data <= f_reg(49);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(50) =>
                        -- NOR R5 R21 R25
                        f_data <= f_reg(50);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(51) =>
                        -- NOP
                        f_data <= f_reg(51);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(52) =>
                        -- SLTIU R6 R19 23581
                        f_data <= f_reg(52);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(53) =>
                        -- SLLV R23 R5 R18
                        f_data <= f_reg(53);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(54) =>
                        -- SLTI R26 R27 29940
                        f_data <= f_reg(54);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(55) =>
                        -- SRL R22 R15 14
                        f_data <= f_reg(55);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(56) =>
                        -- NOP
                        f_data <= f_reg(56);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(57) =>
                        -- SW R19 R0 1096
                        f_data <= f_reg(57);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(58) =>
                        -- ANDI R28 R26 -1792
                        f_data <= f_reg(58);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(59) =>
                        -- NOR R9 R23 R20
                        f_data <= f_reg(59);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(60) =>
                        -- LUI R29 -16537
                        f_data <= f_reg(60);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(61) =>
                        -- SRAV R14 R16 R10
                        f_data <= f_reg(61);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(62) =>
                        -- AND R11 R14 R6
                        f_data <= f_reg(62);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(63) =>
                        -- NOP
                        f_data <= f_reg(63);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(64) =>
                        -- SW R11 R0 1100
                        f_data <= f_reg(64);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(65) =>
                        -- XOR R17 R22 R22
                        f_data <= f_reg(65);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(66) =>
                        -- SW R30 R0 1104
                        f_data <= f_reg(66);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(67) =>
                        -- SLL R12 R0 24
                        f_data <= f_reg(67);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(68) =>
                        -- ADDIU R8 R29 8233
                        f_data <= f_reg(68);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(69) =>
                        -- NOR R4 R17 R24
                        f_data <= f_reg(69);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(70) =>
                        -- SRLV R2 R8 R13
                        f_data <= f_reg(70);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(71) =>
                        -- NOP
                        f_data <= f_reg(71);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(72) =>
                        -- XOR R1 R12 R28
                        f_data <= f_reg(72);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(73) =>
                        -- SLLV R7 R1 R2
                        f_data <= f_reg(73);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(74) =>
                        -- NOP
                        f_data <= f_reg(74);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(75) =>
                        -- SW R9 R0 1108
                        f_data <= f_reg(75);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(76) =>
                        -- SW R7 R0 1112
                        f_data <= f_reg(76);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(77) =>
                        -- SW R4 R0 1116
                        f_data <= f_reg(77);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(78) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(78);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(79) =>
                        -- BGTZ R31 -76
                        f_data <= f_reg(79);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(80) =>
                        -- BEQ R0 R0 454
                        f_data <= f_reg(80);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(81) =>
                        -- LUI R30 999
                        f_data <= f_reg(81);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(82) =>
                        -- LUI R31 999
                        f_data <= f_reg(82);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(83) =>
                        -- SRL R30 R30 16
                        f_data <= f_reg(83);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(84) =>
                        -- SRL R31 R31 16
                        f_data <= f_reg(84);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(85) =>
                        -- LUI R1 -19413
                        f_data <= f_reg(85);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(86) =>
                        -- LUI R15 -19413
                        f_data <= f_reg(86);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(87) =>
                        -- SLTU R2 R1 R0
                        f_data <= f_reg(87);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(88) =>
                        -- SLTU R16 R15 R0
                        f_data <= f_reg(88);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(89) =>
                        -- XORI R3 R2 -14645
                        f_data <= f_reg(89);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(90) =>
                        -- XORI R17 R16 -14645
                        f_data <= f_reg(90);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(91) =>
                        -- SLLV R4 R2 R3
                        f_data <= f_reg(91);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(92) =>
                        -- SLLV R18 R16 R17
                        f_data <= f_reg(92);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(93) =>
                        -- SLT R5 R1 R3
                        f_data <= f_reg(93);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(94) =>
                        -- SLT R19 R15 R17
                        f_data <= f_reg(94);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(95) =>
                        -- SLTIU R6 R4 29340
                        f_data <= f_reg(95);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(96) =>
                        -- SLTIU R20 R18 29340
                        f_data <= f_reg(96);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(97) =>
                        -- SLTIU R7 R6 -11769
                        f_data <= f_reg(97);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(98) =>
                        -- SLTIU R21 R20 -11769
                        f_data <= f_reg(98);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(99) =>
                        -- XOR R8 R7 R7
                        f_data <= f_reg(99);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(100) =>
                        -- XOR R22 R21 R21
                        f_data <= f_reg(100);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(101) =>
                        -- ORI R9 R5 27837
                        f_data <= f_reg(101);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(102) =>
                        -- ORI R23 R19 27837
                        f_data <= f_reg(102);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(103) =>
                        -- SRLV R10 R5 R2
                        f_data <= f_reg(103);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(104) =>
                        -- SRLV R24 R19 R16
                        f_data <= f_reg(104);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(105) =>
                        -- SLL R11 R7 18
                        f_data <= f_reg(105);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(106) =>
                        -- SLL R25 R21 18
                        f_data <= f_reg(106);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(107) =>
                        -- BNE R3 R17 286
                        f_data <= f_reg(107);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(108) =>
                        -- SW R3 R0 1080
                        f_data <= f_reg(108);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(109) =>
                        -- SUB R12 R2 R9
                        f_data <= f_reg(109);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(110) =>
                        -- SUB R26 R16 R23
                        f_data <= f_reg(110);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(111) =>
                        -- OR R13 R4 R0
                        f_data <= f_reg(111);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(112) =>
                        -- OR R27 R18 R0
                        f_data <= f_reg(112);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(113) =>
                        -- ORI R14 R0 30369
                        f_data <= f_reg(113);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(114) =>
                        -- ORI R28 R0 30369
                        f_data <= f_reg(114);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(115) =>
                        -- SLT R1 R12 R13
                        f_data <= f_reg(115);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(116) =>
                        -- SLT R15 R26 R27
                        f_data <= f_reg(116);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(117) =>
                        -- SRLV R12 R1 R8
                        f_data <= f_reg(117);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(118) =>
                        -- SRLV R26 R15 R22
                        f_data <= f_reg(118);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(119) =>
                        -- XOR R8 R2 R1
                        f_data <= f_reg(119);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(120) =>
                        -- XOR R22 R16 R15
                        f_data <= f_reg(120);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(121) =>
                        -- LUI R1 9669
                        f_data <= f_reg(121);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(122) =>
                        -- LUI R15 9669
                        f_data <= f_reg(122);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(123) =>
                        -- BNE R13 R27 270
                        f_data <= f_reg(123);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(124) =>
                        -- SW R13 R0 1120
                        f_data <= f_reg(124);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(125) =>
                        -- SLL R13 R5 21
                        f_data <= f_reg(125);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(126) =>
                        -- SLL R27 R19 21
                        f_data <= f_reg(126);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(127) =>
                        -- BNE R13 R27 266
                        f_data <= f_reg(127);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(128) =>
                        -- SW R13 R0 1124
                        f_data <= f_reg(128);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(129) =>
                        -- LW R13 R0 1120
                        f_data <= f_reg(129);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(130) =>
                        -- LW R27 R0 1120
                        f_data <= f_reg(130);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(131) =>
                        -- BNE R13 R27 -2
                        f_data <= f_reg(131);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(132) =>
                        -- BNE R7 R21 261
                        f_data <= f_reg(132);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(133) =>
                        -- SW R7 R0 1128
                        f_data <= f_reg(133);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(134) =>
                        -- SLTU R7 R13 R14
                        f_data <= f_reg(134);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(135) =>
                        -- SLTU R21 R27 R28
                        f_data <= f_reg(135);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(136) =>
                        -- BNE R13 R27 257
                        f_data <= f_reg(136);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(137) =>
                        -- SW R13 R0 1132
                        f_data <= f_reg(137);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(138) =>
                        -- SUBU R13 R2 R2
                        f_data <= f_reg(138);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(139) =>
                        -- SUBU R27 R16 R16
                        f_data <= f_reg(139);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(140) =>
                        -- SLLV R14 R14 R3
                        f_data <= f_reg(140);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(141) =>
                        -- SLLV R28 R28 R17
                        f_data <= f_reg(141);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(142) =>
                        -- ADDIU R2 R3 -26681
                        f_data <= f_reg(142);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(143) =>
                        -- ADDIU R16 R17 -26681
                        f_data <= f_reg(143);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(144) =>
                        -- SRLV R3 R12 R2
                        f_data <= f_reg(144);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(145) =>
                        -- SRLV R17 R26 R16
                        f_data <= f_reg(145);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(146) =>
                        -- ANDI R12 R7 32377
                        f_data <= f_reg(146);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(147) =>
                        -- ANDI R26 R21 32377
                        f_data <= f_reg(147);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(148) =>
                        -- SUBU R7 R4 R12
                        f_data <= f_reg(148);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(149) =>
                        -- SUBU R21 R18 R26
                        f_data <= f_reg(149);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(150) =>
                        -- BNE R1 R15 243
                        f_data <= f_reg(150);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(151) =>
                        -- SW R1 R0 1084
                        f_data <= f_reg(151);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(152) =>
                        -- SRAV R1 R13 R9
                        f_data <= f_reg(152);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(153) =>
                        -- SRAV R15 R27 R23
                        f_data <= f_reg(153);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(154) =>
                        -- ADDIU R13 R1 -11907
                        f_data <= f_reg(154);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(155) =>
                        -- ADDIU R27 R15 -11907
                        f_data <= f_reg(155);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(156) =>
                        -- BNE R13 R27 237
                        f_data <= f_reg(156);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(157) =>
                        -- SW R13 R0 1136
                        f_data <= f_reg(157);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(158) =>
                        -- OR R13 R12 R10
                        f_data <= f_reg(158);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(159) =>
                        -- OR R27 R26 R24
                        f_data <= f_reg(159);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(160) =>
                        -- ORI R10 R5 27080
                        f_data <= f_reg(160);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(161) =>
                        -- ORI R24 R19 27080
                        f_data <= f_reg(161);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(162) =>
                        -- BNE R13 R27 231
                        f_data <= f_reg(162);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(163) =>
                        -- SW R13 R0 1088
                        f_data <= f_reg(163);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(164) =>
                        -- SRLV R5 R6 R3
                        f_data <= f_reg(164);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(165) =>
                        -- SRLV R19 R20 R17
                        f_data <= f_reg(165);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(166) =>
                        -- OR R6 R1 R2
                        f_data <= f_reg(166);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(167) =>
                        -- OR R20 R15 R16
                        f_data <= f_reg(167);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(168) =>
                        -- BNE R13 R27 225
                        f_data <= f_reg(168);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(169) =>
                        -- SW R13 R0 1092
                        f_data <= f_reg(169);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(170) =>
                        -- ANDI R3 R5 -22366
                        f_data <= f_reg(170);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(171) =>
                        -- ANDI R17 R19 -22366
                        f_data <= f_reg(171);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(172) =>
                        -- SLT R1 R9 R10
                        f_data <= f_reg(172);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(173) =>
                        -- SLT R15 R23 R24
                        f_data <= f_reg(173);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(174) =>
                        -- XOR R4 R3 R4
                        f_data <= f_reg(174);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(175) =>
                        -- XOR R18 R17 R18
                        f_data <= f_reg(175);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(176) =>
                        -- LW R2 R0 1136
                        f_data <= f_reg(176);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(177) =>
                        -- LW R16 R0 1136
                        f_data <= f_reg(177);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(178) =>
                        -- BNE R2 R16 -2
                        f_data <= f_reg(178);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(179) =>
                        -- SLT R13 R14 R2
                        f_data <= f_reg(179);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(180) =>
                        -- SLT R27 R28 R16
                        f_data <= f_reg(180);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(181) =>
                        -- SUBU R9 R11 R8
                        f_data <= f_reg(181);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(182) =>
                        -- SUBU R23 R25 R22
                        f_data <= f_reg(182);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(183) =>
                        -- SRL R10 R3 5
                        f_data <= f_reg(183);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(184) =>
                        -- SRL R24 R17 5
                        f_data <= f_reg(184);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(185) =>
                        -- LW R14 R0 1124
                        f_data <= f_reg(185);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(186) =>
                        -- LW R28 R0 1124
                        f_data <= f_reg(186);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(187) =>
                        -- BNE R14 R28 -2
                        f_data <= f_reg(187);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(188) =>
                        -- SUB R11 R1 R14
                        f_data <= f_reg(188);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(189) =>
                        -- SUB R25 R15 R28
                        f_data <= f_reg(189);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(190) =>
                        -- LW R8 R0 1128
                        f_data <= f_reg(190);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(191) =>
                        -- LW R22 R0 1128
                        f_data <= f_reg(191);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(192) =>
                        -- BNE R8 R22 -2
                        f_data <= f_reg(192);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(193) =>
                        -- XOR R3 R4 R8
                        f_data <= f_reg(193);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(194) =>
                        -- XOR R17 R18 R22
                        f_data <= f_reg(194);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(195) =>
                        -- LW R1 R0 1132
                        f_data <= f_reg(195);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(196) =>
                        -- LW R15 R0 1132
                        f_data <= f_reg(196);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(197) =>
                        -- BNE R1 R15 -2
                        f_data <= f_reg(197);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(198) =>
                        -- ADDU R4 R9 R1
                        f_data <= f_reg(198);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(199) =>
                        -- ADDU R18 R23 R15
                        f_data <= f_reg(199);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(200) =>
                        -- SLLV R9 R6 R8
                        f_data <= f_reg(200);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(201) =>
                        -- SLLV R23 R20 R22
                        f_data <= f_reg(201);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(202) =>
                        -- SLTIU R6 R10 25015
                        f_data <= f_reg(202);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(203) =>
                        -- SLTIU R20 R24 25015
                        f_data <= f_reg(203);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(204) =>
                        -- NOR R8 R9 R7
                        f_data <= f_reg(204);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(205) =>
                        -- NOR R22 R23 R21
                        f_data <= f_reg(205);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(206) =>
                        -- NOP
                        f_data <= f_reg(206);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(207) =>
                        -- NOP
                        f_data <= f_reg(207);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(208) =>
                        -- SLTIU R10 R14 23581
                        f_data <= f_reg(208);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(209) =>
                        -- SLTIU R24 R28 23581
                        f_data <= f_reg(209);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(210) =>
                        -- SLLV R9 R8 R4
                        f_data <= f_reg(210);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(211) =>
                        -- SLLV R23 R22 R18
                        f_data <= f_reg(211);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(212) =>
                        -- SLTI R7 R2 29940
                        f_data <= f_reg(212);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(213) =>
                        -- SLTI R21 R16 29940
                        f_data <= f_reg(213);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(214) =>
                        -- SRL R8 R13 14
                        f_data <= f_reg(214);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(215) =>
                        -- SRL R22 R27 14
                        f_data <= f_reg(215);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(216) =>
                        -- NOP
                        f_data <= f_reg(216);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(217) =>
                        -- NOP
                        f_data <= f_reg(217);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(218) =>
                        -- BNE R14 R28 175
                        f_data <= f_reg(218);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(219) =>
                        -- SW R14 R0 1096
                        f_data <= f_reg(219);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(220) =>
                        -- ANDI R4 R7 -1792
                        f_data <= f_reg(220);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(221) =>
                        -- ANDI R18 R21 -1792
                        f_data <= f_reg(221);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(222) =>
                        -- NOR R2 R9 R3
                        f_data <= f_reg(222);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(223) =>
                        -- NOR R16 R23 R17
                        f_data <= f_reg(223);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(224) =>
                        -- LUI R13 -16537
                        f_data <= f_reg(224);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(225) =>
                        -- LUI R27 -16537
                        f_data <= f_reg(225);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(226) =>
                        -- SRAV R14 R11 R6
                        f_data <= f_reg(226);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(227) =>
                        -- SRAV R28 R25 R20
                        f_data <= f_reg(227);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(228) =>
                        -- AND R7 R14 R10
                        f_data <= f_reg(228);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(229) =>
                        -- AND R21 R28 R24
                        f_data <= f_reg(229);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(230) =>
                        -- NOP
                        f_data <= f_reg(230);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(231) =>
                        -- NOP
                        f_data <= f_reg(231);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(232) =>
                        -- BNE R7 R21 161
                        f_data <= f_reg(232);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(233) =>
                        -- SW R7 R0 1100
                        f_data <= f_reg(233);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(234) =>
                        -- XOR R9 R8 R8
                        f_data <= f_reg(234);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(235) =>
                        -- XOR R23 R22 R22
                        f_data <= f_reg(235);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(236) =>
                        -- BNE R5 R19 157
                        f_data <= f_reg(236);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(237) =>
                        -- SW R5 R0 1104
                        f_data <= f_reg(237);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(238) =>
                        -- SLL R3 R0 24
                        f_data <= f_reg(238);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(239) =>
                        -- SLL R17 R0 24
                        f_data <= f_reg(239);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(240) =>
                        -- ADDIU R11 R13 8233
                        f_data <= f_reg(240);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(241) =>
                        -- ADDIU R25 R27 8233
                        f_data <= f_reg(241);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(242) =>
                        -- NOR R6 R9 R12
                        f_data <= f_reg(242);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(243) =>
                        -- NOR R20 R23 R26
                        f_data <= f_reg(243);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(244) =>
                        -- SRLV R14 R11 R1
                        f_data <= f_reg(244);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(245) =>
                        -- SRLV R28 R25 R15
                        f_data <= f_reg(245);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(246) =>
                        -- NOP
                        f_data <= f_reg(246);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(247) =>
                        -- NOP
                        f_data <= f_reg(247);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(248) =>
                        -- XOR R10 R3 R4
                        f_data <= f_reg(248);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(249) =>
                        -- XOR R24 R17 R18
                        f_data <= f_reg(249);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(250) =>
                        -- SLLV R7 R10 R14
                        f_data <= f_reg(250);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(251) =>
                        -- SLLV R21 R24 R28
                        f_data <= f_reg(251);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(252) =>
                        -- NOP
                        f_data <= f_reg(252);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(253) =>
                        -- NOP
                        f_data <= f_reg(253);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(254) =>
                        -- BNE R2 R16 139
                        f_data <= f_reg(254);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(255) =>
                        -- SW R2 R0 1108
                        f_data <= f_reg(255);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(256) =>
                        -- BNE R7 R21 137
                        f_data <= f_reg(256);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(257) =>
                        -- SW R7 R0 1112
                        f_data <= f_reg(257);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(258) =>
                        -- BNE R6 R20 135
                        f_data <= f_reg(258);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(259) =>
                        -- SW R6 R0 1116
                        f_data <= f_reg(259);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(260) =>
                        -- ADDI R29 R30 -250
                        f_data <= f_reg(260);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(261) =>
                        -- BEQ R29 R0 25
                        f_data <= f_reg(261);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(262) =>
                        -- ADDI R29 R30 -500
                        f_data <= f_reg(262);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(263) =>
                        -- BEQ R29 R0 23
                        f_data <= f_reg(263);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(264) =>
                        -- ADDI R29 R30 -750
                        f_data <= f_reg(264);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(265) =>
                        -- BEQ R29 R0 21
                        f_data <= f_reg(265);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(266) =>
                        -- ADDI R30 R30 -1
                        f_data <= f_reg(266);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(267) =>
                        -- ADDI R31 R31 -1
                        f_data <= f_reg(267);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(268) =>
                        -- BNE R30 R31 125
                        f_data <= f_reg(268);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(269) =>
                        -- BGTZ R31 -184
                        f_data <= f_reg(269);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(270) =>
                        -- BEQ R0 R0 264
                        f_data <= f_reg(270);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(271) =>
                        -- NOP
                        f_data <= f_reg(271);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(272) =>
                        -- NOP
                        f_data <= f_reg(272);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(273) =>
                        -- NOP
                        f_data <= f_reg(273);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(274) =>
                        -- NOP
                        f_data <= f_reg(274);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(275) =>
                        -- NOP
                        f_data <= f_reg(275);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(276) =>
                        -- NOP
                        f_data <= f_reg(276);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(277) =>
                        -- NOP
                        f_data <= f_reg(277);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(278) =>
                        -- NOP
                        f_data <= f_reg(278);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(279) =>
                        -- NOP
                        f_data <= f_reg(279);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(280) =>
                        -- NOP
                        f_data <= f_reg(280);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(281) =>
                        -- NOP
                        f_data <= f_reg(281);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(282) =>
                        -- NOP
                        f_data <= f_reg(282);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(283) =>
                        -- NOP
                        f_data <= f_reg(283);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(284) =>
                        -- NOP
                        f_data <= f_reg(284);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(285) =>
                        -- NOP
                        f_data <= f_reg(285);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(286) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(286);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(287) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(287);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(288) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(288);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(289) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(289);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(290) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(290);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(291) =>
                        -- BNE R1 R15 102
                        f_data <= f_reg(291);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(292) =>
                        -- SW R1 R29 1872
                        f_data <= f_reg(292);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(293) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(293);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(294) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(294);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(295) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(295);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(296) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(296);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(297) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(297);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(298) =>
                        -- BNE R2 R16 95
                        f_data <= f_reg(298);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(299) =>
                        -- SW R2 R29 1876
                        f_data <= f_reg(299);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(300) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(300);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(301) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(301);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(302) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(302);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(303) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(303);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(304) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(304);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(305) =>
                        -- BNE R3 R17 88
                        f_data <= f_reg(305);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(306) =>
                        -- SW R3 R29 1880
                        f_data <= f_reg(306);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(307) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(307);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(308) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(308);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(309) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(309);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(310) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(310);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(311) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(311);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(312) =>
                        -- BNE R4 R18 81
                        f_data <= f_reg(312);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(313) =>
                        -- SW R4 R29 1884
                        f_data <= f_reg(313);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(314) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(314);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(315) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(315);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(316) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(316);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(317) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(317);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(318) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(318);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(319) =>
                        -- BNE R5 R19 74
                        f_data <= f_reg(319);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(320) =>
                        -- SW R5 R29 1888
                        f_data <= f_reg(320);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(321) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(321);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(322) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(322);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(323) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(323);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(324) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(324);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(325) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(325);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(326) =>
                        -- BNE R6 R20 67
                        f_data <= f_reg(326);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(327) =>
                        -- SW R6 R29 1892
                        f_data <= f_reg(327);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(328) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(328);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(329) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(329);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(330) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(330);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(331) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(331);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(332) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(332);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(333) =>
                        -- BNE R7 R21 60
                        f_data <= f_reg(333);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(334) =>
                        -- SW R7 R29 1896
                        f_data <= f_reg(334);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(335) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(335);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(336) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(336);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(337) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(337);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(338) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(338);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(339) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(339);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(340) =>
                        -- BNE R8 R22 53
                        f_data <= f_reg(340);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(341) =>
                        -- SW R8 R29 1900
                        f_data <= f_reg(341);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(342) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(342);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(343) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(343);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(344) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(344);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(345) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(345);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(346) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(346);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(347) =>
                        -- BNE R9 R23 46
                        f_data <= f_reg(347);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(348) =>
                        -- SW R9 R29 1904
                        f_data <= f_reg(348);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(349) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(349);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(350) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(350);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(351) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(351);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(352) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(352);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(353) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(353);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(354) =>
                        -- BNE R10 R24 39
                        f_data <= f_reg(354);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(355) =>
                        -- SW R10 R29 1908
                        f_data <= f_reg(355);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(356) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(356);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(357) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(357);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(358) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(358);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(359) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(359);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(360) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(360);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(361) =>
                        -- BNE R11 R25 32
                        f_data <= f_reg(361);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(362) =>
                        -- SW R11 R29 1912
                        f_data <= f_reg(362);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(363) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(363);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(364) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(364);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(365) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(365);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(366) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(366);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(367) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(367);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(368) =>
                        -- BNE R12 R26 25
                        f_data <= f_reg(368);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(369) =>
                        -- SW R12 R29 1916
                        f_data <= f_reg(369);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(370) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(370);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(371) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(371);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(372) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(372);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(373) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(373);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(374) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(374);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(375) =>
                        -- BNE R13 R27 18
                        f_data <= f_reg(375);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(376) =>
                        -- SW R13 R29 1920
                        f_data <= f_reg(376);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(377) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(377);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(378) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(378);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(379) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(379);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(380) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(380);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(381) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(381);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(382) =>
                        -- BNE R14 R28 11
                        f_data <= f_reg(382);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(383) =>
                        -- SW R14 R29 1924
                        f_data <= f_reg(383);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(384) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(384);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(385) =>
                        -- BGTZ R29 3
                        f_data <= f_reg(385);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(386) =>
                        -- ADDI R29 R0 60
                        f_data <= f_reg(386);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(387) =>
                        -- BEQ R0 R0 2
                        f_data <= f_reg(387);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(388) =>
                        -- ADDI R29 R0 0
                        f_data <= f_reg(388);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(389) =>
                        -- BNE R30 R31 4
                        f_data <= f_reg(389);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(390) =>
                        -- SW R30 R29 1928
                        f_data <= f_reg(390);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(391) =>
                        -- SW R29 R0 1992
                        f_data <= f_reg(391);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(392) =>
                        -- BEQ R0 R0 -126
                        f_data <= f_reg(392);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(393) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(393);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(394) =>
                        -- LW R1 R29 1872
                        f_data <= f_reg(394);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(395) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(395);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(396) =>
                        -- LW R15 R29 1872
                        f_data <= f_reg(396);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(397) =>
                        -- BNE R1 R15 -4
                        f_data <= f_reg(397);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(398) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(398);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(399) =>
                        -- LW R2 R29 1876
                        f_data <= f_reg(399);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(400) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(400);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(401) =>
                        -- LW R16 R29 1876
                        f_data <= f_reg(401);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(402) =>
                        -- BNE R2 R16 -4
                        f_data <= f_reg(402);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(403) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(403);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(404) =>
                        -- LW R3 R29 1880
                        f_data <= f_reg(404);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(405) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(405);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(406) =>
                        -- LW R17 R29 1880
                        f_data <= f_reg(406);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(407) =>
                        -- BNE R3 R17 -4
                        f_data <= f_reg(407);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(408) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(408);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(409) =>
                        -- LW R4 R29 1884
                        f_data <= f_reg(409);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(410) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(410);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(411) =>
                        -- LW R18 R29 1884
                        f_data <= f_reg(411);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(412) =>
                        -- BNE R4 R18 -4
                        f_data <= f_reg(412);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(413) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(413);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(414) =>
                        -- LW R5 R29 1888
                        f_data <= f_reg(414);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(415) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(415);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(416) =>
                        -- LW R19 R29 1888
                        f_data <= f_reg(416);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(417) =>
                        -- BNE R5 R19 -4
                        f_data <= f_reg(417);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(418) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(418);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(419) =>
                        -- LW R6 R29 1892
                        f_data <= f_reg(419);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(420) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(420);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(421) =>
                        -- LW R20 R29 1892
                        f_data <= f_reg(421);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(422) =>
                        -- BNE R6 R20 -4
                        f_data <= f_reg(422);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(423) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(423);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(424) =>
                        -- LW R7 R29 1896
                        f_data <= f_reg(424);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(425) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(425);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(426) =>
                        -- LW R21 R29 1896
                        f_data <= f_reg(426);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(427) =>
                        -- BNE R7 R21 -4
                        f_data <= f_reg(427);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(428) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(428);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(429) =>
                        -- LW R8 R29 1900
                        f_data <= f_reg(429);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(430) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(430);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(431) =>
                        -- LW R22 R29 1900
                        f_data <= f_reg(431);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(432) =>
                        -- BNE R8 R22 -4
                        f_data <= f_reg(432);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(433) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(433);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(434) =>
                        -- LW R9 R29 1904
                        f_data <= f_reg(434);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(435) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(435);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(436) =>
                        -- LW R23 R29 1904
                        f_data <= f_reg(436);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(437) =>
                        -- BNE R9 R23 -4
                        f_data <= f_reg(437);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(438) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(438);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(439) =>
                        -- LW R10 R29 1908
                        f_data <= f_reg(439);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(440) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(440);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(441) =>
                        -- LW R24 R29 1908
                        f_data <= f_reg(441);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(442) =>
                        -- BNE R10 R24 -4
                        f_data <= f_reg(442);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(443) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(443);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(444) =>
                        -- LW R11 R29 1912
                        f_data <= f_reg(444);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(445) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(445);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(446) =>
                        -- LW R25 R29 1912
                        f_data <= f_reg(446);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(447) =>
                        -- BNE R11 R25 -4
                        f_data <= f_reg(447);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(448) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(448);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(449) =>
                        -- LW R12 R29 1916
                        f_data <= f_reg(449);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(450) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(450);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(451) =>
                        -- LW R26 R29 1916
                        f_data <= f_reg(451);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(452) =>
                        -- BNE R12 R26 -4
                        f_data <= f_reg(452);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(453) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(453);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(454) =>
                        -- LW R13 R29 1920
                        f_data <= f_reg(454);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(455) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(455);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(456) =>
                        -- LW R27 R29 1920
                        f_data <= f_reg(456);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(457) =>
                        -- BNE R13 R27 -4
                        f_data <= f_reg(457);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(458) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(458);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(459) =>
                        -- LW R14 R29 1924
                        f_data <= f_reg(459);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(460) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(460);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(461) =>
                        -- LW R28 R29 1924
                        f_data <= f_reg(461);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(462) =>
                        -- BNE R14 R28 -4
                        f_data <= f_reg(462);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(463) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(463);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(464) =>
                        -- LW R30 R29 1928
                        f_data <= f_reg(464);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(465) =>
                        -- LW R29 R0 1992
                        f_data <= f_reg(465);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(466) =>
                        -- LW R31 R29 1928
                        f_data <= f_reg(466);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(467) =>
                        -- BNE R30 R31 -4
                        f_data <= f_reg(467);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(468) =>
                        -- BEQ R0 R0 -202
                        f_data <= f_reg(468);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(469) =>
                        -- NOP
                        f_data <= f_reg(469);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(470) =>
                        -- NOP
                        f_data <= f_reg(470);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(471) =>
                        -- NOP
                        f_data <= f_reg(471);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(472) =>
                        -- NOP
                        f_data <= f_reg(472);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(473) =>
                        -- NOP
                        f_data <= f_reg(473);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(474) =>
                        -- NOP
                        f_data <= f_reg(474);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(475) =>
                        -- NOP
                        f_data <= f_reg(475);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(476) =>
                        -- NOP
                        f_data <= f_reg(476);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(477) =>
                        -- NOP
                        f_data <= f_reg(477);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(478) =>
                        -- NOP
                        f_data <= f_reg(478);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(479) =>
                        -- NOP
                        f_data <= f_reg(479);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(480) =>
                        -- NOP
                        f_data <= f_reg(480);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(481) =>
                        -- NOP
                        f_data <= f_reg(481);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(482) =>
                        -- NOP
                        f_data <= f_reg(482);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(483) =>
                        -- NOP
                        f_data <= f_reg(483);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(484) =>
                        -- NOP
                        f_data <= f_reg(484);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(485) =>
                        -- NOP
                        f_data <= f_reg(485);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(486) =>
                        -- NOP
                        f_data <= f_reg(486);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(487) =>
                        -- NOP
                        f_data <= f_reg(487);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(488) =>
                        -- NOP
                        f_data <= f_reg(488);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(489) =>
                        -- NOP
                        f_data <= f_reg(489);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(490) =>
                        -- NOP
                        f_data <= f_reg(490);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(491) =>
                        -- NOP
                        f_data <= f_reg(491);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(492) =>
                        -- NOP
                        f_data <= f_reg(492);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(493) =>
                        -- NOP
                        f_data <= f_reg(493);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(494) =>
                        -- NOP
                        f_data <= f_reg(494);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(495) =>
                        -- NOP
                        f_data <= f_reg(495);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(496) =>
                        -- NOP
                        f_data <= f_reg(496);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(497) =>
                        -- NOP
                        f_data <= f_reg(497);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(498) =>
                        -- NOP
                        f_data <= f_reg(498);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(499) =>
                        -- NOP
                        f_data <= f_reg(499);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(500) =>
                        -- NOP
                        f_data <= f_reg(500);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(501) =>
                        -- NOP
                        f_data <= f_reg(501);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(502) =>
                        -- NOP
                        f_data <= f_reg(502);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(503) =>
                        -- NOP
                        f_data <= f_reg(503);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(504) =>
                        -- NOP
                        f_data <= f_reg(504);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(505) =>
                        -- NOP
                        f_data <= f_reg(505);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(506) =>
                        -- NOP
                        f_data <= f_reg(506);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(507) =>
                        -- NOP
                        f_data <= f_reg(507);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(508) =>
                        -- NOP
                        f_data <= f_reg(508);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(509) =>
                        -- NOP
                        f_data <= f_reg(509);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(510) =>
                        -- NOP
                        f_data <= f_reg(510);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(511) =>
                        -- NOP
                        f_data <= f_reg(511);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(512) =>
                        -- NOP
                        f_data <= f_reg(512);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(513) =>
                        -- NOP
                        f_data <= f_reg(513);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(514) =>
                        -- NOP
                        f_data <= f_reg(514);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(515) =>
                        -- NOP
                        f_data <= f_reg(515);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(516) =>
                        -- NOP
                        f_data <= f_reg(516);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(517) =>
                        -- NOP
                        f_data <= f_reg(517);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(518) =>
                        -- NOP
                        f_data <= f_reg(518);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(519) =>
                        -- NOP
                        f_data <= f_reg(519);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(520) =>
                        -- NOP
                        f_data <= f_reg(520);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(521) =>
                        -- NOP
                        f_data <= f_reg(521);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(522) =>
                        -- NOP
                        f_data <= f_reg(522);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(523) =>
                        -- NOP
                        f_data <= f_reg(523);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(524) =>
                        -- NOP
                        f_data <= f_reg(524);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(525) =>
                        -- NOP
                        f_data <= f_reg(525);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(526) =>
                        -- NOP
                        f_data <= f_reg(526);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(527) =>
                        -- NOP
                        f_data <= f_reg(527);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(528) =>
                        -- NOP
                        f_data <= f_reg(528);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(529) =>
                        -- NOP
                        f_data <= f_reg(529);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(530) =>
                        -- NOP
                        f_data <= f_reg(530);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(531) =>
                        -- NOP
                        f_data <= f_reg(531);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(532) =>
                        -- NOP
                        f_data <= f_reg(532);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(533) =>
                        -- NOP
                        f_data <= f_reg(533);
                        f_MEM_READY <= '1';
                        f_DONE <= '0';
                     when k_prog(534) =>
                        -- End of Program
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011011010000101011";
                        f_reg(4) <= "00000000001000000001000000101011";
                        f_reg(5) <= "00111000010000111100011011001011";
                        f_reg(6) <= "00000000011000100010000000000100";
                        f_reg(7) <= "00000000001000110010100000101010";
                        f_reg(8) <= "00101100100001100111001010011100";
                        f_reg(9) <= "00101100110001111101001000000111";
                        f_reg(10) <= "00000000111001110100000000100110";
                        f_reg(11) <= "00110100101010010110110010111101";
                        f_reg(12) <= "00000000010001010101000000000110";
                        f_reg(13) <= "00000000000001110101110010000000";
                        f_reg(14) <= "10101100000000110000010000111000";
                        f_reg(15) <= "00000000010010010110000000100010";
                        f_reg(16) <= "00000000100000000110100000100101";
                        f_reg(17) <= "00110100000011100111011010100001";
                        f_reg(18) <= "00000001100011010111100000101010";
                        f_reg(19) <= "00000001000011111000000000000110";
                        f_reg(20) <= "00000000010011111000100000100110";
                        f_reg(21) <= "00111100000100100010010111000101";
                        f_reg(22) <= "00000000000001011001110101000000";
                        f_reg(23) <= "00000001101011101010000000101011";
                        f_reg(24) <= "00000000010000101010100000100011";
                        f_reg(25) <= "00000000011011100111000000000100";
                        f_reg(26) <= "00100100011101101001011111000111";
                        f_reg(27) <= "00000010110100001011100000000110";
                        f_reg(28) <= "00110010100110000111111001111001";
                        f_reg(29) <= "00000000100110001100100000100011";
                        f_reg(30) <= "10101100000100100000010000111100";
                        f_reg(31) <= "00000001001101011101000000000111";
                        f_reg(32) <= "00100111010110111101000101111101";
                        f_reg(33) <= "00000011000010101110000000100101";
                        f_reg(34) <= "00110100101111010110100111001000";
                        f_reg(35) <= "10101100000111000000010001000000";
                        f_reg(36) <= "00000010111001101111000000000110";
                        f_reg(37) <= "00000011010101100000100000100101";
                        f_reg(38) <= "10101100000111000000010001000100";
                        f_reg(39) <= "00110011110011001010100010100010";
                        f_reg(40) <= "00000001001111010100000000101010";
                        f_reg(41) <= "00000001100001000010000000100110";
                        f_reg(42) <= "00000001110110110111100000101010";
                        f_reg(43) <= "00000001011100010001000000100011";
                        f_reg(44) <= "00000000000011000001100101000010";
                        f_reg(45) <= "00000001000100111000000000100010";
                        f_reg(46) <= "00000000100001111010000000100110";
                        f_reg(47) <= "00000000010011011001000000100001";
                        f_reg(48) <= "00000000111000011010100000000100";
                        f_reg(49) <= "00101100011010100110000110110111";
                        f_reg(50) <= "00000010101110010010100000100111";
                        f_reg(51) <= "00000000000000000000000000000000";
                        f_reg(52) <= "00101110011001100101110000011101";
                        f_reg(53) <= "00000010010001011011100000000100";
                        f_reg(54) <= "00101011011110100111010011110100";
                        f_reg(55) <= "00000000000011111011001110000010";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "10101100000100110000010001001000";
                        f_reg(58) <= "00110011010111001111100100000000";
                        f_reg(59) <= "00000010111101000100100000100111";
                        f_reg(60) <= "00111100000111011011111101100111";
                        f_reg(61) <= "00000001010100000111000000000111";
                        f_reg(62) <= "00000001110001100101100000100100";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000010110000010001001100";
                        f_reg(65) <= "00000010110101101000100000100110";
                        f_reg(66) <= "10101100000111100000010001010000";
                        f_reg(67) <= "00000000000000000110011000000000";
                        f_reg(68) <= "00100111101010000010000000101001";
                        f_reg(69) <= "00000010001110000010000000100111";
                        f_reg(70) <= "00000001101010000001000000000110";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000001100111000000100000100110";
                        f_reg(73) <= "00000000010000010011100000000100";
                        f_reg(74) <= "00000000000000000000000000000000";
                        f_reg(75) <= "10101100000010010000010001010100";
                        f_reg(76) <= "10101100000001110000010001011000";
                        f_reg(77) <= "10101100000001000000010001011100";
                        f_reg(78) <= "00100011111111111111111111111111";
                        f_reg(79) <= "00011111111000001111111110110100";
                        f_reg(80) <= "00010000000000000000000111000110";
                        f_reg(81) <= "00111100000111100000001111100111";
                        f_reg(82) <= "00111100000111110000001111100111";
                        f_reg(83) <= "00000000000111101111010000000010";
                        f_reg(84) <= "00000000000111111111110000000010";
                        f_reg(85) <= "00111100000000011011010000101011";
                        f_reg(86) <= "00111100000011111011010000101011";
                        f_reg(87) <= "00000000001000000001000000101011";
                        f_reg(88) <= "00000001111000001000000000101011";
                        f_reg(89) <= "00111000010000111100011011001011";
                        f_reg(90) <= "00111010000100011100011011001011";
                        f_reg(91) <= "00000000011000100010000000000100";
                        f_reg(92) <= "00000010001100001001000000000100";
                        f_reg(93) <= "00000000001000110010100000101010";
                        f_reg(94) <= "00000001111100011001100000101010";
                        f_reg(95) <= "00101100100001100111001010011100";
                        f_reg(96) <= "00101110010101000111001010011100";
                        f_reg(97) <= "00101100110001111101001000000111";
                        f_reg(98) <= "00101110100101011101001000000111";
                        f_reg(99) <= "00000000111001110100000000100110";
                        f_reg(100) <= "00000010101101011011000000100110";
                        f_reg(101) <= "00110100101010010110110010111101";
                        f_reg(102) <= "00110110011101110110110010111101";
                        f_reg(103) <= "00000000010001010101000000000110";
                        f_reg(104) <= "00000010000100111100000000000110";
                        f_reg(105) <= "00000000000001110101110010000000";
                        f_reg(106) <= "00000000000101011100110010000000";
                        f_reg(107) <= "00010100011100010000000100011110";
                        f_reg(108) <= "10101100000000110000010000111000";
                        f_reg(109) <= "00000000010010010110000000100010";
                        f_reg(110) <= "00000010000101111101000000100010";
                        f_reg(111) <= "00000000100000000110100000100101";
                        f_reg(112) <= "00000010010000001101100000100101";
                        f_reg(113) <= "00110100000011100111011010100001";
                        f_reg(114) <= "00110100000111000111011010100001";
                        f_reg(115) <= "00000001100011010000100000101010";
                        f_reg(116) <= "00000011010110110111100000101010";
                        f_reg(117) <= "00000001000000010110000000000110";
                        f_reg(118) <= "00000010110011111101000000000110";
                        f_reg(119) <= "00000000010000010100000000100110";
                        f_reg(120) <= "00000010000011111011000000100110";
                        f_reg(121) <= "00111100000000010010010111000101";
                        f_reg(122) <= "00111100000011110010010111000101";
                        f_reg(123) <= "00010101101110110000000100001110";
                        f_reg(124) <= "10101100000011010000010001100000";
                        f_reg(125) <= "00000000000001010110110101000000";
                        f_reg(126) <= "00000000000100111101110101000000";
                        f_reg(127) <= "00010101101110110000000100001010";
                        f_reg(128) <= "10101100000011010000010001100100";
                        f_reg(129) <= "10001100000011010000010001100000";
                        f_reg(130) <= "10001100000110110000010001100000";
                        f_reg(131) <= "00010101101110111111111111111110";
                        f_reg(132) <= "00010100111101010000000100000101";
                        f_reg(133) <= "10101100000001110000010001101000";
                        f_reg(134) <= "00000001101011100011100000101011";
                        f_reg(135) <= "00000011011111001010100000101011";
                        f_reg(136) <= "00010101101110110000000100000001";
                        f_reg(137) <= "10101100000011010000010001101100";
                        f_reg(138) <= "00000000010000100110100000100011";
                        f_reg(139) <= "00000010000100001101100000100011";
                        f_reg(140) <= "00000000011011100111000000000100";
                        f_reg(141) <= "00000010001111001110000000000100";
                        f_reg(142) <= "00100100011000101001011111000111";
                        f_reg(143) <= "00100110001100001001011111000111";
                        f_reg(144) <= "00000000010011000001100000000110";
                        f_reg(145) <= "00000010000110101000100000000110";
                        f_reg(146) <= "00110000111011000111111001111001";
                        f_reg(147) <= "00110010101110100111111001111001";
                        f_reg(148) <= "00000000100011000011100000100011";
                        f_reg(149) <= "00000010010110101010100000100011";
                        f_reg(150) <= "00010100001011110000000011110011";
                        f_reg(151) <= "10101100000000010000010000111100";
                        f_reg(152) <= "00000001001011010000100000000111";
                        f_reg(153) <= "00000010111110110111100000000111";
                        f_reg(154) <= "00100100001011011101000101111101";
                        f_reg(155) <= "00100101111110111101000101111101";
                        f_reg(156) <= "00010101101110110000000011101101";
                        f_reg(157) <= "10101100000011010000010001110000";
                        f_reg(158) <= "00000001100010100110100000100101";
                        f_reg(159) <= "00000011010110001101100000100101";
                        f_reg(160) <= "00110100101010100110100111001000";
                        f_reg(161) <= "00110110011110000110100111001000";
                        f_reg(162) <= "00010101101110110000000011100111";
                        f_reg(163) <= "10101100000011010000010001000000";
                        f_reg(164) <= "00000000011001100010100000000110";
                        f_reg(165) <= "00000010001101001001100000000110";
                        f_reg(166) <= "00000000001000100011000000100101";
                        f_reg(167) <= "00000001111100001010000000100101";
                        f_reg(168) <= "00010101101110110000000011100001";
                        f_reg(169) <= "10101100000011010000010001000100";
                        f_reg(170) <= "00110000101000111010100010100010";
                        f_reg(171) <= "00110010011100011010100010100010";
                        f_reg(172) <= "00000001001010100000100000101010";
                        f_reg(173) <= "00000010111110000111100000101010";
                        f_reg(174) <= "00000000011001000010000000100110";
                        f_reg(175) <= "00000010001100101001000000100110";
                        f_reg(176) <= "10001100000000100000010001110000";
                        f_reg(177) <= "10001100000100000000010001110000";
                        f_reg(178) <= "00010100010100001111111111111110";
                        f_reg(179) <= "00000001110000100110100000101010";
                        f_reg(180) <= "00000011100100001101100000101010";
                        f_reg(181) <= "00000001011010000100100000100011";
                        f_reg(182) <= "00000011001101101011100000100011";
                        f_reg(183) <= "00000000000000110101000101000010";
                        f_reg(184) <= "00000000000100011100000101000010";
                        f_reg(185) <= "10001100000011100000010001100100";
                        f_reg(186) <= "10001100000111000000010001100100";
                        f_reg(187) <= "00010101110111001111111111111110";
                        f_reg(188) <= "00000000001011100101100000100010";
                        f_reg(189) <= "00000001111111001100100000100010";
                        f_reg(190) <= "10001100000010000000010001101000";
                        f_reg(191) <= "10001100000101100000010001101000";
                        f_reg(192) <= "00010101000101101111111111111110";
                        f_reg(193) <= "00000000100010000001100000100110";
                        f_reg(194) <= "00000010010101101000100000100110";
                        f_reg(195) <= "10001100000000010000010001101100";
                        f_reg(196) <= "10001100000011110000010001101100";
                        f_reg(197) <= "00010100001011111111111111111110";
                        f_reg(198) <= "00000001001000010010000000100001";
                        f_reg(199) <= "00000010111011111001000000100001";
                        f_reg(200) <= "00000001000001100100100000000100";
                        f_reg(201) <= "00000010110101001011100000000100";
                        f_reg(202) <= "00101101010001100110000110110111";
                        f_reg(203) <= "00101111000101000110000110110111";
                        f_reg(204) <= "00000001001001110100000000100111";
                        f_reg(205) <= "00000010111101011011000000100111";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101101110010100101110000011101";
                        f_reg(209) <= "00101111100110000101110000011101";
                        f_reg(210) <= "00000000100010000100100000000100";
                        f_reg(211) <= "00000010010101101011100000000100";
                        f_reg(212) <= "00101000010001110111010011110100";
                        f_reg(213) <= "00101010000101010111010011110100";
                        f_reg(214) <= "00000000000011010100001110000010";
                        f_reg(215) <= "00000000000110111011001110000010";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "00010101110111000000000010101111";
                        f_reg(219) <= "10101100000011100000010001001000";
                        f_reg(220) <= "00110000111001001111100100000000";
                        f_reg(221) <= "00110010101100101111100100000000";
                        f_reg(222) <= "00000001001000110001000000100111";
                        f_reg(223) <= "00000010111100011000000000100111";
                        f_reg(224) <= "00111100000011011011111101100111";
                        f_reg(225) <= "00111100000110111011111101100111";
                        f_reg(226) <= "00000000110010110111000000000111";
                        f_reg(227) <= "00000010100110011110000000000111";
                        f_reg(228) <= "00000001110010100011100000100100";
                        f_reg(229) <= "00000011100110001010100000100100";
                        f_reg(230) <= "00000000000000000000000000000000";
                        f_reg(231) <= "00000000000000000000000000000000";
                        f_reg(232) <= "00010100111101010000000010100001";
                        f_reg(233) <= "10101100000001110000010001001100";
                        f_reg(234) <= "00000001000010000100100000100110";
                        f_reg(235) <= "00000010110101101011100000100110";
                        f_reg(236) <= "00010100101100110000000010011101";
                        f_reg(237) <= "10101100000001010000010001010000";
                        f_reg(238) <= "00000000000000000001111000000000";
                        f_reg(239) <= "00000000000000001000111000000000";
                        f_reg(240) <= "00100101101010110010000000101001";
                        f_reg(241) <= "00100111011110010010000000101001";
                        f_reg(242) <= "00000001001011000011000000100111";
                        f_reg(243) <= "00000010111110101010000000100111";
                        f_reg(244) <= "00000000001010110111000000000110";
                        f_reg(245) <= "00000001111110011110000000000110";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00000000011001000101000000100110";
                        f_reg(249) <= "00000010001100101100000000100110";
                        f_reg(250) <= "00000001110010100011100000000100";
                        f_reg(251) <= "00000011100110001010100000000100";
                        f_reg(252) <= "00000000000000000000000000000000";
                        f_reg(253) <= "00000000000000000000000000000000";
                        f_reg(254) <= "00010100010100000000000010001011";
                        f_reg(255) <= "10101100000000100000010001010100";
                        f_reg(256) <= "00010100111101010000000010001001";
                        f_reg(257) <= "10101100000001110000010001011000";
                        f_reg(258) <= "00010100110101000000000010000111";
                        f_reg(259) <= "10101100000001100000010001011100";
                        f_reg(260) <= "00100011110111011111111100000110";
                        f_reg(261) <= "00010011101000000000000000011001";
                        f_reg(262) <= "00100011110111011111111000001100";
                        f_reg(263) <= "00010011101000000000000000010111";
                        f_reg(264) <= "00100011110111011111110100010010";
                        f_reg(265) <= "00010011101000000000000000010101";
                        f_reg(266) <= "00100011110111101111111111111111";
                        f_reg(267) <= "00100011111111111111111111111111";
                        f_reg(268) <= "00010111110111110000000001111101";
                        f_reg(269) <= "00011111111000001111111101001000";
                        f_reg(270) <= "00010000000000000000000100001000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "10001100000111010000011111001000";
                        f_reg(287) <= "00011111101000000000000000000011";
                        f_reg(288) <= "00100000000111010000000000111100";
                        f_reg(289) <= "00010000000000000000000000000010";
                        f_reg(290) <= "00100000000111010000000000000000";
                        f_reg(291) <= "00010100001011110000000001100110";
                        f_reg(292) <= "10101111101000010000011101010000";
                        f_reg(293) <= "10001100000111010000011111001000";
                        f_reg(294) <= "00011111101000000000000000000011";
                        f_reg(295) <= "00100000000111010000000000111100";
                        f_reg(296) <= "00010000000000000000000000000010";
                        f_reg(297) <= "00100000000111010000000000000000";
                        f_reg(298) <= "00010100010100000000000001011111";
                        f_reg(299) <= "10101111101000100000011101010100";
                        f_reg(300) <= "10001100000111010000011111001000";
                        f_reg(301) <= "00011111101000000000000000000011";
                        f_reg(302) <= "00100000000111010000000000111100";
                        f_reg(303) <= "00010000000000000000000000000010";
                        f_reg(304) <= "00100000000111010000000000000000";
                        f_reg(305) <= "00010100011100010000000001011000";
                        f_reg(306) <= "10101111101000110000011101011000";
                        f_reg(307) <= "10001100000111010000011111001000";
                        f_reg(308) <= "00011111101000000000000000000011";
                        f_reg(309) <= "00100000000111010000000000111100";
                        f_reg(310) <= "00010000000000000000000000000010";
                        f_reg(311) <= "00100000000111010000000000000000";
                        f_reg(312) <= "00010100100100100000000001010001";
                        f_reg(313) <= "10101111101001000000011101011100";
                        f_reg(314) <= "10001100000111010000011111001000";
                        f_reg(315) <= "00011111101000000000000000000011";
                        f_reg(316) <= "00100000000111010000000000111100";
                        f_reg(317) <= "00010000000000000000000000000010";
                        f_reg(318) <= "00100000000111010000000000000000";
                        f_reg(319) <= "00010100101100110000000001001010";
                        f_reg(320) <= "10101111101001010000011101100000";
                        f_reg(321) <= "10001100000111010000011111001000";
                        f_reg(322) <= "00011111101000000000000000000011";
                        f_reg(323) <= "00100000000111010000000000111100";
                        f_reg(324) <= "00010000000000000000000000000010";
                        f_reg(325) <= "00100000000111010000000000000000";
                        f_reg(326) <= "00010100110101000000000001000011";
                        f_reg(327) <= "10101111101001100000011101100100";
                        f_reg(328) <= "10001100000111010000011111001000";
                        f_reg(329) <= "00011111101000000000000000000011";
                        f_reg(330) <= "00100000000111010000000000111100";
                        f_reg(331) <= "00010000000000000000000000000010";
                        f_reg(332) <= "00100000000111010000000000000000";
                        f_reg(333) <= "00010100111101010000000000111100";
                        f_reg(334) <= "10101111101001110000011101101000";
                        f_reg(335) <= "10001100000111010000011111001000";
                        f_reg(336) <= "00011111101000000000000000000011";
                        f_reg(337) <= "00100000000111010000000000111100";
                        f_reg(338) <= "00010000000000000000000000000010";
                        f_reg(339) <= "00100000000111010000000000000000";
                        f_reg(340) <= "00010101000101100000000000110101";
                        f_reg(341) <= "10101111101010000000011101101100";
                        f_reg(342) <= "10001100000111010000011111001000";
                        f_reg(343) <= "00011111101000000000000000000011";
                        f_reg(344) <= "00100000000111010000000000111100";
                        f_reg(345) <= "00010000000000000000000000000010";
                        f_reg(346) <= "00100000000111010000000000000000";
                        f_reg(347) <= "00010101001101110000000000101110";
                        f_reg(348) <= "10101111101010010000011101110000";
                        f_reg(349) <= "10001100000111010000011111001000";
                        f_reg(350) <= "00011111101000000000000000000011";
                        f_reg(351) <= "00100000000111010000000000111100";
                        f_reg(352) <= "00010000000000000000000000000010";
                        f_reg(353) <= "00100000000111010000000000000000";
                        f_reg(354) <= "00010101010110000000000000100111";
                        f_reg(355) <= "10101111101010100000011101110100";
                        f_reg(356) <= "10001100000111010000011111001000";
                        f_reg(357) <= "00011111101000000000000000000011";
                        f_reg(358) <= "00100000000111010000000000111100";
                        f_reg(359) <= "00010000000000000000000000000010";
                        f_reg(360) <= "00100000000111010000000000000000";
                        f_reg(361) <= "00010101011110010000000000100000";
                        f_reg(362) <= "10101111101010110000011101111000";
                        f_reg(363) <= "10001100000111010000011111001000";
                        f_reg(364) <= "00011111101000000000000000000011";
                        f_reg(365) <= "00100000000111010000000000111100";
                        f_reg(366) <= "00010000000000000000000000000010";
                        f_reg(367) <= "00100000000111010000000000000000";
                        f_reg(368) <= "00010101100110100000000000011001";
                        f_reg(369) <= "10101111101011000000011101111100";
                        f_reg(370) <= "10001100000111010000011111001000";
                        f_reg(371) <= "00011111101000000000000000000011";
                        f_reg(372) <= "00100000000111010000000000111100";
                        f_reg(373) <= "00010000000000000000000000000010";
                        f_reg(374) <= "00100000000111010000000000000000";
                        f_reg(375) <= "00010101101110110000000000010010";
                        f_reg(376) <= "10101111101011010000011110000000";
                        f_reg(377) <= "10001100000111010000011111001000";
                        f_reg(378) <= "00011111101000000000000000000011";
                        f_reg(379) <= "00100000000111010000000000111100";
                        f_reg(380) <= "00010000000000000000000000000010";
                        f_reg(381) <= "00100000000111010000000000000000";
                        f_reg(382) <= "00010101110111000000000000001011";
                        f_reg(383) <= "10101111101011100000011110000100";
                        f_reg(384) <= "10001100000111010000011111001000";
                        f_reg(385) <= "00011111101000000000000000000011";
                        f_reg(386) <= "00100000000111010000000000111100";
                        f_reg(387) <= "00010000000000000000000000000010";
                        f_reg(388) <= "00100000000111010000000000000000";
                        f_reg(389) <= "00010111110111110000000000000100";
                        f_reg(390) <= "10101111101111100000011110001000";
                        f_reg(391) <= "10101100000111010000011111001000";
                        f_reg(392) <= "00010000000000001111111110000010";
                        f_reg(393) <= "10001100000111010000011111001000";
                        f_reg(394) <= "10001111101000010000011101010000";
                        f_reg(395) <= "10001100000111010000011111001000";
                        f_reg(396) <= "10001111101011110000011101010000";
                        f_reg(397) <= "00010100001011111111111111111100";
                        f_reg(398) <= "10001100000111010000011111001000";
                        f_reg(399) <= "10001111101000100000011101010100";
                        f_reg(400) <= "10001100000111010000011111001000";
                        f_reg(401) <= "10001111101100000000011101010100";
                        f_reg(402) <= "00010100010100001111111111111100";
                        f_reg(403) <= "10001100000111010000011111001000";
                        f_reg(404) <= "10001111101000110000011101011000";
                        f_reg(405) <= "10001100000111010000011111001000";
                        f_reg(406) <= "10001111101100010000011101011000";
                        f_reg(407) <= "00010100011100011111111111111100";
                        f_reg(408) <= "10001100000111010000011111001000";
                        f_reg(409) <= "10001111101001000000011101011100";
                        f_reg(410) <= "10001100000111010000011111001000";
                        f_reg(411) <= "10001111101100100000011101011100";
                        f_reg(412) <= "00010100100100101111111111111100";
                        f_reg(413) <= "10001100000111010000011111001000";
                        f_reg(414) <= "10001111101001010000011101100000";
                        f_reg(415) <= "10001100000111010000011111001000";
                        f_reg(416) <= "10001111101100110000011101100000";
                        f_reg(417) <= "00010100101100111111111111111100";
                        f_reg(418) <= "10001100000111010000011111001000";
                        f_reg(419) <= "10001111101001100000011101100100";
                        f_reg(420) <= "10001100000111010000011111001000";
                        f_reg(421) <= "10001111101101000000011101100100";
                        f_reg(422) <= "00010100110101001111111111111100";
                        f_reg(423) <= "10001100000111010000011111001000";
                        f_reg(424) <= "10001111101001110000011101101000";
                        f_reg(425) <= "10001100000111010000011111001000";
                        f_reg(426) <= "10001111101101010000011101101000";
                        f_reg(427) <= "00010100111101011111111111111100";
                        f_reg(428) <= "10001100000111010000011111001000";
                        f_reg(429) <= "10001111101010000000011101101100";
                        f_reg(430) <= "10001100000111010000011111001000";
                        f_reg(431) <= "10001111101101100000011101101100";
                        f_reg(432) <= "00010101000101101111111111111100";
                        f_reg(433) <= "10001100000111010000011111001000";
                        f_reg(434) <= "10001111101010010000011101110000";
                        f_reg(435) <= "10001100000111010000011111001000";
                        f_reg(436) <= "10001111101101110000011101110000";
                        f_reg(437) <= "00010101001101111111111111111100";
                        f_reg(438) <= "10001100000111010000011111001000";
                        f_reg(439) <= "10001111101010100000011101110100";
                        f_reg(440) <= "10001100000111010000011111001000";
                        f_reg(441) <= "10001111101110000000011101110100";
                        f_reg(442) <= "00010101010110001111111111111100";
                        f_reg(443) <= "10001100000111010000011111001000";
                        f_reg(444) <= "10001111101010110000011101111000";
                        f_reg(445) <= "10001100000111010000011111001000";
                        f_reg(446) <= "10001111101110010000011101111000";
                        f_reg(447) <= "00010101011110011111111111111100";
                        f_reg(448) <= "10001100000111010000011111001000";
                        f_reg(449) <= "10001111101011000000011101111100";
                        f_reg(450) <= "10001100000111010000011111001000";
                        f_reg(451) <= "10001111101110100000011101111100";
                        f_reg(452) <= "00010101100110101111111111111100";
                        f_reg(453) <= "10001100000111010000011111001000";
                        f_reg(454) <= "10001111101011010000011110000000";
                        f_reg(455) <= "10001100000111010000011111001000";
                        f_reg(456) <= "10001111101110110000011110000000";
                        f_reg(457) <= "00010101101110111111111111111100";
                        f_reg(458) <= "10001100000111010000011111001000";
                        f_reg(459) <= "10001111101011100000011110000100";
                        f_reg(460) <= "10001100000111010000011111001000";
                        f_reg(461) <= "10001111101111000000011110000100";
                        f_reg(462) <= "00010101110111001111111111111100";
                        f_reg(463) <= "10001100000111010000011111001000";
                        f_reg(464) <= "10001111101111100000011110001000";
                        f_reg(465) <= "10001100000111010000011111001000";
                        f_reg(466) <= "10001111101111110000011110001000";
                        f_reg(467) <= "00010111110111111111111111111100";
                        f_reg(468) <= "00010000000000001111111100110110";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000001111100111";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                     when others =>
                        -- Jump to Location Outside of Program -- An error has occured
                        f_data <= B"00000000000000000000000000000000";
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_timeout_flag <= '0';
                        f_recovery_flag <= '0';
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011011010000101011";
                        f_reg(4) <= "00000000001000000001000000101011";
                        f_reg(5) <= "00111000010000111100011011001011";
                        f_reg(6) <= "00000000011000100010000000000100";
                        f_reg(7) <= "00000000001000110010100000101010";
                        f_reg(8) <= "00101100100001100111001010011100";
                        f_reg(9) <= "00101100110001111101001000000111";
                        f_reg(10) <= "00000000111001110100000000100110";
                        f_reg(11) <= "00110100101010010110110010111101";
                        f_reg(12) <= "00000000010001010101000000000110";
                        f_reg(13) <= "00000000000001110101110010000000";
                        f_reg(14) <= "10101100000000110000010000111000";
                        f_reg(15) <= "00000000010010010110000000100010";
                        f_reg(16) <= "00000000100000000110100000100101";
                        f_reg(17) <= "00110100000011100111011010100001";
                        f_reg(18) <= "00000001100011010111100000101010";
                        f_reg(19) <= "00000001000011111000000000000110";
                        f_reg(20) <= "00000000010011111000100000100110";
                        f_reg(21) <= "00111100000100100010010111000101";
                        f_reg(22) <= "00000000000001011001110101000000";
                        f_reg(23) <= "00000001101011101010000000101011";
                        f_reg(24) <= "00000000010000101010100000100011";
                        f_reg(25) <= "00000000011011100111000000000100";
                        f_reg(26) <= "00100100011101101001011111000111";
                        f_reg(27) <= "00000010110100001011100000000110";
                        f_reg(28) <= "00110010100110000111111001111001";
                        f_reg(29) <= "00000000100110001100100000100011";
                        f_reg(30) <= "10101100000100100000010000111100";
                        f_reg(31) <= "00000001001101011101000000000111";
                        f_reg(32) <= "00100111010110111101000101111101";
                        f_reg(33) <= "00000011000010101110000000100101";
                        f_reg(34) <= "00110100101111010110100111001000";
                        f_reg(35) <= "10101100000111000000010001000000";
                        f_reg(36) <= "00000010111001101111000000000110";
                        f_reg(37) <= "00000011010101100000100000100101";
                        f_reg(38) <= "10101100000111000000010001000100";
                        f_reg(39) <= "00110011110011001010100010100010";
                        f_reg(40) <= "00000001001111010100000000101010";
                        f_reg(41) <= "00000001100001000010000000100110";
                        f_reg(42) <= "00000001110110110111100000101010";
                        f_reg(43) <= "00000001011100010001000000100011";
                        f_reg(44) <= "00000000000011000001100101000010";
                        f_reg(45) <= "00000001000100111000000000100010";
                        f_reg(46) <= "00000000100001111010000000100110";
                        f_reg(47) <= "00000000010011011001000000100001";
                        f_reg(48) <= "00000000111000011010100000000100";
                        f_reg(49) <= "00101100011010100110000110110111";
                        f_reg(50) <= "00000010101110010010100000100111";
                        f_reg(51) <= "00000000000000000000000000000000";
                        f_reg(52) <= "00101110011001100101110000011101";
                        f_reg(53) <= "00000010010001011011100000000100";
                        f_reg(54) <= "00101011011110100111010011110100";
                        f_reg(55) <= "00000000000011111011001110000010";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "10101100000100110000010001001000";
                        f_reg(58) <= "00110011010111001111100100000000";
                        f_reg(59) <= "00000010111101000100100000100111";
                        f_reg(60) <= "00111100000111011011111101100111";
                        f_reg(61) <= "00000001010100000111000000000111";
                        f_reg(62) <= "00000001110001100101100000100100";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000010110000010001001100";
                        f_reg(65) <= "00000010110101101000100000100110";
                        f_reg(66) <= "10101100000111100000010001010000";
                        f_reg(67) <= "00000000000000000110011000000000";
                        f_reg(68) <= "00100111101010000010000000101001";
                        f_reg(69) <= "00000010001110000010000000100111";
                        f_reg(70) <= "00000001101010000001000000000110";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000001100111000000100000100110";
                        f_reg(73) <= "00000000010000010011100000000100";
                        f_reg(74) <= "00000000000000000000000000000000";
                        f_reg(75) <= "10101100000010010000010001010100";
                        f_reg(76) <= "10101100000001110000010001011000";
                        f_reg(77) <= "10101100000001000000010001011100";
                        f_reg(78) <= "00100011111111111111111111111111";
                        f_reg(79) <= "00011111111000001111111110110100";
                        f_reg(80) <= "00010000000000000000000111000110";
                        f_reg(81) <= "00111100000111100000001111100111";
                        f_reg(82) <= "00111100000111110000001111100111";
                        f_reg(83) <= "00000000000111101111010000000010";
                        f_reg(84) <= "00000000000111111111110000000010";
                        f_reg(85) <= "00111100000000011011010000101011";
                        f_reg(86) <= "00111100000011111011010000101011";
                        f_reg(87) <= "00000000001000000001000000101011";
                        f_reg(88) <= "00000001111000001000000000101011";
                        f_reg(89) <= "00111000010000111100011011001011";
                        f_reg(90) <= "00111010000100011100011011001011";
                        f_reg(91) <= "00000000011000100010000000000100";
                        f_reg(92) <= "00000010001100001001000000000100";
                        f_reg(93) <= "00000000001000110010100000101010";
                        f_reg(94) <= "00000001111100011001100000101010";
                        f_reg(95) <= "00101100100001100111001010011100";
                        f_reg(96) <= "00101110010101000111001010011100";
                        f_reg(97) <= "00101100110001111101001000000111";
                        f_reg(98) <= "00101110100101011101001000000111";
                        f_reg(99) <= "00000000111001110100000000100110";
                        f_reg(100) <= "00000010101101011011000000100110";
                        f_reg(101) <= "00110100101010010110110010111101";
                        f_reg(102) <= "00110110011101110110110010111101";
                        f_reg(103) <= "00000000010001010101000000000110";
                        f_reg(104) <= "00000010000100111100000000000110";
                        f_reg(105) <= "00000000000001110101110010000000";
                        f_reg(106) <= "00000000000101011100110010000000";
                        f_reg(107) <= "00010100011100010000000100011110";
                        f_reg(108) <= "10101100000000110000010000111000";
                        f_reg(109) <= "00000000010010010110000000100010";
                        f_reg(110) <= "00000010000101111101000000100010";
                        f_reg(111) <= "00000000100000000110100000100101";
                        f_reg(112) <= "00000010010000001101100000100101";
                        f_reg(113) <= "00110100000011100111011010100001";
                        f_reg(114) <= "00110100000111000111011010100001";
                        f_reg(115) <= "00000001100011010000100000101010";
                        f_reg(116) <= "00000011010110110111100000101010";
                        f_reg(117) <= "00000001000000010110000000000110";
                        f_reg(118) <= "00000010110011111101000000000110";
                        f_reg(119) <= "00000000010000010100000000100110";
                        f_reg(120) <= "00000010000011111011000000100110";
                        f_reg(121) <= "00111100000000010010010111000101";
                        f_reg(122) <= "00111100000011110010010111000101";
                        f_reg(123) <= "00010101101110110000000100001110";
                        f_reg(124) <= "10101100000011010000010001100000";
                        f_reg(125) <= "00000000000001010110110101000000";
                        f_reg(126) <= "00000000000100111101110101000000";
                        f_reg(127) <= "00010101101110110000000100001010";
                        f_reg(128) <= "10101100000011010000010001100100";
                        f_reg(129) <= "10001100000011010000010001100000";
                        f_reg(130) <= "10001100000110110000010001100000";
                        f_reg(131) <= "00010101101110111111111111111110";
                        f_reg(132) <= "00010100111101010000000100000101";
                        f_reg(133) <= "10101100000001110000010001101000";
                        f_reg(134) <= "00000001101011100011100000101011";
                        f_reg(135) <= "00000011011111001010100000101011";
                        f_reg(136) <= "00010101101110110000000100000001";
                        f_reg(137) <= "10101100000011010000010001101100";
                        f_reg(138) <= "00000000010000100110100000100011";
                        f_reg(139) <= "00000010000100001101100000100011";
                        f_reg(140) <= "00000000011011100111000000000100";
                        f_reg(141) <= "00000010001111001110000000000100";
                        f_reg(142) <= "00100100011000101001011111000111";
                        f_reg(143) <= "00100110001100001001011111000111";
                        f_reg(144) <= "00000000010011000001100000000110";
                        f_reg(145) <= "00000010000110101000100000000110";
                        f_reg(146) <= "00110000111011000111111001111001";
                        f_reg(147) <= "00110010101110100111111001111001";
                        f_reg(148) <= "00000000100011000011100000100011";
                        f_reg(149) <= "00000010010110101010100000100011";
                        f_reg(150) <= "00010100001011110000000011110011";
                        f_reg(151) <= "10101100000000010000010000111100";
                        f_reg(152) <= "00000001001011010000100000000111";
                        f_reg(153) <= "00000010111110110111100000000111";
                        f_reg(154) <= "00100100001011011101000101111101";
                        f_reg(155) <= "00100101111110111101000101111101";
                        f_reg(156) <= "00010101101110110000000011101101";
                        f_reg(157) <= "10101100000011010000010001110000";
                        f_reg(158) <= "00000001100010100110100000100101";
                        f_reg(159) <= "00000011010110001101100000100101";
                        f_reg(160) <= "00110100101010100110100111001000";
                        f_reg(161) <= "00110110011110000110100111001000";
                        f_reg(162) <= "00010101101110110000000011100111";
                        f_reg(163) <= "10101100000011010000010001000000";
                        f_reg(164) <= "00000000011001100010100000000110";
                        f_reg(165) <= "00000010001101001001100000000110";
                        f_reg(166) <= "00000000001000100011000000100101";
                        f_reg(167) <= "00000001111100001010000000100101";
                        f_reg(168) <= "00010101101110110000000011100001";
                        f_reg(169) <= "10101100000011010000010001000100";
                        f_reg(170) <= "00110000101000111010100010100010";
                        f_reg(171) <= "00110010011100011010100010100010";
                        f_reg(172) <= "00000001001010100000100000101010";
                        f_reg(173) <= "00000010111110000111100000101010";
                        f_reg(174) <= "00000000011001000010000000100110";
                        f_reg(175) <= "00000010001100101001000000100110";
                        f_reg(176) <= "10001100000000100000010001110000";
                        f_reg(177) <= "10001100000100000000010001110000";
                        f_reg(178) <= "00010100010100001111111111111110";
                        f_reg(179) <= "00000001110000100110100000101010";
                        f_reg(180) <= "00000011100100001101100000101010";
                        f_reg(181) <= "00000001011010000100100000100011";
                        f_reg(182) <= "00000011001101101011100000100011";
                        f_reg(183) <= "00000000000000110101000101000010";
                        f_reg(184) <= "00000000000100011100000101000010";
                        f_reg(185) <= "10001100000011100000010001100100";
                        f_reg(186) <= "10001100000111000000010001100100";
                        f_reg(187) <= "00010101110111001111111111111110";
                        f_reg(188) <= "00000000001011100101100000100010";
                        f_reg(189) <= "00000001111111001100100000100010";
                        f_reg(190) <= "10001100000010000000010001101000";
                        f_reg(191) <= "10001100000101100000010001101000";
                        f_reg(192) <= "00010101000101101111111111111110";
                        f_reg(193) <= "00000000100010000001100000100110";
                        f_reg(194) <= "00000010010101101000100000100110";
                        f_reg(195) <= "10001100000000010000010001101100";
                        f_reg(196) <= "10001100000011110000010001101100";
                        f_reg(197) <= "00010100001011111111111111111110";
                        f_reg(198) <= "00000001001000010010000000100001";
                        f_reg(199) <= "00000010111011111001000000100001";
                        f_reg(200) <= "00000001000001100100100000000100";
                        f_reg(201) <= "00000010110101001011100000000100";
                        f_reg(202) <= "00101101010001100110000110110111";
                        f_reg(203) <= "00101111000101000110000110110111";
                        f_reg(204) <= "00000001001001110100000000100111";
                        f_reg(205) <= "00000010111101011011000000100111";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101101110010100101110000011101";
                        f_reg(209) <= "00101111100110000101110000011101";
                        f_reg(210) <= "00000000100010000100100000000100";
                        f_reg(211) <= "00000010010101101011100000000100";
                        f_reg(212) <= "00101000010001110111010011110100";
                        f_reg(213) <= "00101010000101010111010011110100";
                        f_reg(214) <= "00000000000011010100001110000010";
                        f_reg(215) <= "00000000000110111011001110000010";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "00010101110111000000000010101111";
                        f_reg(219) <= "10101100000011100000010001001000";
                        f_reg(220) <= "00110000111001001111100100000000";
                        f_reg(221) <= "00110010101100101111100100000000";
                        f_reg(222) <= "00000001001000110001000000100111";
                        f_reg(223) <= "00000010111100011000000000100111";
                        f_reg(224) <= "00111100000011011011111101100111";
                        f_reg(225) <= "00111100000110111011111101100111";
                        f_reg(226) <= "00000000110010110111000000000111";
                        f_reg(227) <= "00000010100110011110000000000111";
                        f_reg(228) <= "00000001110010100011100000100100";
                        f_reg(229) <= "00000011100110001010100000100100";
                        f_reg(230) <= "00000000000000000000000000000000";
                        f_reg(231) <= "00000000000000000000000000000000";
                        f_reg(232) <= "00010100111101010000000010100001";
                        f_reg(233) <= "10101100000001110000010001001100";
                        f_reg(234) <= "00000001000010000100100000100110";
                        f_reg(235) <= "00000010110101101011100000100110";
                        f_reg(236) <= "00010100101100110000000010011101";
                        f_reg(237) <= "10101100000001010000010001010000";
                        f_reg(238) <= "00000000000000000001111000000000";
                        f_reg(239) <= "00000000000000001000111000000000";
                        f_reg(240) <= "00100101101010110010000000101001";
                        f_reg(241) <= "00100111011110010010000000101001";
                        f_reg(242) <= "00000001001011000011000000100111";
                        f_reg(243) <= "00000010111110101010000000100111";
                        f_reg(244) <= "00000000001010110111000000000110";
                        f_reg(245) <= "00000001111110011110000000000110";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00000000011001000101000000100110";
                        f_reg(249) <= "00000010001100101100000000100110";
                        f_reg(250) <= "00000001110010100011100000000100";
                        f_reg(251) <= "00000011100110001010100000000100";
                        f_reg(252) <= "00000000000000000000000000000000";
                        f_reg(253) <= "00000000000000000000000000000000";
                        f_reg(254) <= "00010100010100000000000010001011";
                        f_reg(255) <= "10101100000000100000010001010100";
                        f_reg(256) <= "00010100111101010000000010001001";
                        f_reg(257) <= "10101100000001110000010001011000";
                        f_reg(258) <= "00010100110101000000000010000111";
                        f_reg(259) <= "10101100000001100000010001011100";
                        f_reg(260) <= "00100011110111011111111100000110";
                        f_reg(261) <= "00010011101000000000000000011001";
                        f_reg(262) <= "00100011110111011111111000001100";
                        f_reg(263) <= "00010011101000000000000000010111";
                        f_reg(264) <= "00100011110111011111110100010010";
                        f_reg(265) <= "00010011101000000000000000010101";
                        f_reg(266) <= "00100011110111101111111111111111";
                        f_reg(267) <= "00100011111111111111111111111111";
                        f_reg(268) <= "00010111110111110000000001111101";
                        f_reg(269) <= "00011111111000001111111101001000";
                        f_reg(270) <= "00010000000000000000000100001000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "10001100000111010000011111001000";
                        f_reg(287) <= "00011111101000000000000000000011";
                        f_reg(288) <= "00100000000111010000000000111100";
                        f_reg(289) <= "00010000000000000000000000000010";
                        f_reg(290) <= "00100000000111010000000000000000";
                        f_reg(291) <= "00010100001011110000000001100110";
                        f_reg(292) <= "10101111101000010000011101010000";
                        f_reg(293) <= "10001100000111010000011111001000";
                        f_reg(294) <= "00011111101000000000000000000011";
                        f_reg(295) <= "00100000000111010000000000111100";
                        f_reg(296) <= "00010000000000000000000000000010";
                        f_reg(297) <= "00100000000111010000000000000000";
                        f_reg(298) <= "00010100010100000000000001011111";
                        f_reg(299) <= "10101111101000100000011101010100";
                        f_reg(300) <= "10001100000111010000011111001000";
                        f_reg(301) <= "00011111101000000000000000000011";
                        f_reg(302) <= "00100000000111010000000000111100";
                        f_reg(303) <= "00010000000000000000000000000010";
                        f_reg(304) <= "00100000000111010000000000000000";
                        f_reg(305) <= "00010100011100010000000001011000";
                        f_reg(306) <= "10101111101000110000011101011000";
                        f_reg(307) <= "10001100000111010000011111001000";
                        f_reg(308) <= "00011111101000000000000000000011";
                        f_reg(309) <= "00100000000111010000000000111100";
                        f_reg(310) <= "00010000000000000000000000000010";
                        f_reg(311) <= "00100000000111010000000000000000";
                        f_reg(312) <= "00010100100100100000000001010001";
                        f_reg(313) <= "10101111101001000000011101011100";
                        f_reg(314) <= "10001100000111010000011111001000";
                        f_reg(315) <= "00011111101000000000000000000011";
                        f_reg(316) <= "00100000000111010000000000111100";
                        f_reg(317) <= "00010000000000000000000000000010";
                        f_reg(318) <= "00100000000111010000000000000000";
                        f_reg(319) <= "00010100101100110000000001001010";
                        f_reg(320) <= "10101111101001010000011101100000";
                        f_reg(321) <= "10001100000111010000011111001000";
                        f_reg(322) <= "00011111101000000000000000000011";
                        f_reg(323) <= "00100000000111010000000000111100";
                        f_reg(324) <= "00010000000000000000000000000010";
                        f_reg(325) <= "00100000000111010000000000000000";
                        f_reg(326) <= "00010100110101000000000001000011";
                        f_reg(327) <= "10101111101001100000011101100100";
                        f_reg(328) <= "10001100000111010000011111001000";
                        f_reg(329) <= "00011111101000000000000000000011";
                        f_reg(330) <= "00100000000111010000000000111100";
                        f_reg(331) <= "00010000000000000000000000000010";
                        f_reg(332) <= "00100000000111010000000000000000";
                        f_reg(333) <= "00010100111101010000000000111100";
                        f_reg(334) <= "10101111101001110000011101101000";
                        f_reg(335) <= "10001100000111010000011111001000";
                        f_reg(336) <= "00011111101000000000000000000011";
                        f_reg(337) <= "00100000000111010000000000111100";
                        f_reg(338) <= "00010000000000000000000000000010";
                        f_reg(339) <= "00100000000111010000000000000000";
                        f_reg(340) <= "00010101000101100000000000110101";
                        f_reg(341) <= "10101111101010000000011101101100";
                        f_reg(342) <= "10001100000111010000011111001000";
                        f_reg(343) <= "00011111101000000000000000000011";
                        f_reg(344) <= "00100000000111010000000000111100";
                        f_reg(345) <= "00010000000000000000000000000010";
                        f_reg(346) <= "00100000000111010000000000000000";
                        f_reg(347) <= "00010101001101110000000000101110";
                        f_reg(348) <= "10101111101010010000011101110000";
                        f_reg(349) <= "10001100000111010000011111001000";
                        f_reg(350) <= "00011111101000000000000000000011";
                        f_reg(351) <= "00100000000111010000000000111100";
                        f_reg(352) <= "00010000000000000000000000000010";
                        f_reg(353) <= "00100000000111010000000000000000";
                        f_reg(354) <= "00010101010110000000000000100111";
                        f_reg(355) <= "10101111101010100000011101110100";
                        f_reg(356) <= "10001100000111010000011111001000";
                        f_reg(357) <= "00011111101000000000000000000011";
                        f_reg(358) <= "00100000000111010000000000111100";
                        f_reg(359) <= "00010000000000000000000000000010";
                        f_reg(360) <= "00100000000111010000000000000000";
                        f_reg(361) <= "00010101011110010000000000100000";
                        f_reg(362) <= "10101111101010110000011101111000";
                        f_reg(363) <= "10001100000111010000011111001000";
                        f_reg(364) <= "00011111101000000000000000000011";
                        f_reg(365) <= "00100000000111010000000000111100";
                        f_reg(366) <= "00010000000000000000000000000010";
                        f_reg(367) <= "00100000000111010000000000000000";
                        f_reg(368) <= "00010101100110100000000000011001";
                        f_reg(369) <= "10101111101011000000011101111100";
                        f_reg(370) <= "10001100000111010000011111001000";
                        f_reg(371) <= "00011111101000000000000000000011";
                        f_reg(372) <= "00100000000111010000000000111100";
                        f_reg(373) <= "00010000000000000000000000000010";
                        f_reg(374) <= "00100000000111010000000000000000";
                        f_reg(375) <= "00010101101110110000000000010010";
                        f_reg(376) <= "10101111101011010000011110000000";
                        f_reg(377) <= "10001100000111010000011111001000";
                        f_reg(378) <= "00011111101000000000000000000011";
                        f_reg(379) <= "00100000000111010000000000111100";
                        f_reg(380) <= "00010000000000000000000000000010";
                        f_reg(381) <= "00100000000111010000000000000000";
                        f_reg(382) <= "00010101110111000000000000001011";
                        f_reg(383) <= "10101111101011100000011110000100";
                        f_reg(384) <= "10001100000111010000011111001000";
                        f_reg(385) <= "00011111101000000000000000000011";
                        f_reg(386) <= "00100000000111010000000000111100";
                        f_reg(387) <= "00010000000000000000000000000010";
                        f_reg(388) <= "00100000000111010000000000000000";
                        f_reg(389) <= "00010111110111110000000000000100";
                        f_reg(390) <= "10101111101111100000011110001000";
                        f_reg(391) <= "10101100000111010000011111001000";
                        f_reg(392) <= "00010000000000001111111110000010";
                        f_reg(393) <= "10001100000111010000011111001000";
                        f_reg(394) <= "10001111101000010000011101010000";
                        f_reg(395) <= "10001100000111010000011111001000";
                        f_reg(396) <= "10001111101011110000011101010000";
                        f_reg(397) <= "00010100001011111111111111111100";
                        f_reg(398) <= "10001100000111010000011111001000";
                        f_reg(399) <= "10001111101000100000011101010100";
                        f_reg(400) <= "10001100000111010000011111001000";
                        f_reg(401) <= "10001111101100000000011101010100";
                        f_reg(402) <= "00010100010100001111111111111100";
                        f_reg(403) <= "10001100000111010000011111001000";
                        f_reg(404) <= "10001111101000110000011101011000";
                        f_reg(405) <= "10001100000111010000011111001000";
                        f_reg(406) <= "10001111101100010000011101011000";
                        f_reg(407) <= "00010100011100011111111111111100";
                        f_reg(408) <= "10001100000111010000011111001000";
                        f_reg(409) <= "10001111101001000000011101011100";
                        f_reg(410) <= "10001100000111010000011111001000";
                        f_reg(411) <= "10001111101100100000011101011100";
                        f_reg(412) <= "00010100100100101111111111111100";
                        f_reg(413) <= "10001100000111010000011111001000";
                        f_reg(414) <= "10001111101001010000011101100000";
                        f_reg(415) <= "10001100000111010000011111001000";
                        f_reg(416) <= "10001111101100110000011101100000";
                        f_reg(417) <= "00010100101100111111111111111100";
                        f_reg(418) <= "10001100000111010000011111001000";
                        f_reg(419) <= "10001111101001100000011101100100";
                        f_reg(420) <= "10001100000111010000011111001000";
                        f_reg(421) <= "10001111101101000000011101100100";
                        f_reg(422) <= "00010100110101001111111111111100";
                        f_reg(423) <= "10001100000111010000011111001000";
                        f_reg(424) <= "10001111101001110000011101101000";
                        f_reg(425) <= "10001100000111010000011111001000";
                        f_reg(426) <= "10001111101101010000011101101000";
                        f_reg(427) <= "00010100111101011111111111111100";
                        f_reg(428) <= "10001100000111010000011111001000";
                        f_reg(429) <= "10001111101010000000011101101100";
                        f_reg(430) <= "10001100000111010000011111001000";
                        f_reg(431) <= "10001111101101100000011101101100";
                        f_reg(432) <= "00010101000101101111111111111100";
                        f_reg(433) <= "10001100000111010000011111001000";
                        f_reg(434) <= "10001111101010010000011101110000";
                        f_reg(435) <= "10001100000111010000011111001000";
                        f_reg(436) <= "10001111101101110000011101110000";
                        f_reg(437) <= "00010101001101111111111111111100";
                        f_reg(438) <= "10001100000111010000011111001000";
                        f_reg(439) <= "10001111101010100000011101110100";
                        f_reg(440) <= "10001100000111010000011111001000";
                        f_reg(441) <= "10001111101110000000011101110100";
                        f_reg(442) <= "00010101010110001111111111111100";
                        f_reg(443) <= "10001100000111010000011111001000";
                        f_reg(444) <= "10001111101010110000011101111000";
                        f_reg(445) <= "10001100000111010000011111001000";
                        f_reg(446) <= "10001111101110010000011101111000";
                        f_reg(447) <= "00010101011110011111111111111100";
                        f_reg(448) <= "10001100000111010000011111001000";
                        f_reg(449) <= "10001111101011000000011101111100";
                        f_reg(450) <= "10001100000111010000011111001000";
                        f_reg(451) <= "10001111101110100000011101111100";
                        f_reg(452) <= "00010101100110101111111111111100";
                        f_reg(453) <= "10001100000111010000011111001000";
                        f_reg(454) <= "10001111101011010000011110000000";
                        f_reg(455) <= "10001100000111010000011111001000";
                        f_reg(456) <= "10001111101110110000011110000000";
                        f_reg(457) <= "00010101101110111111111111111100";
                        f_reg(458) <= "10001100000111010000011111001000";
                        f_reg(459) <= "10001111101011100000011110000100";
                        f_reg(460) <= "10001100000111010000011111001000";
                        f_reg(461) <= "10001111101111000000011110000100";
                        f_reg(462) <= "00010101110111001111111111111100";
                        f_reg(463) <= "10001100000111010000011111001000";
                        f_reg(464) <= "10001111101111100000011110001000";
                        f_reg(465) <= "10001100000111010000011111001000";
                        f_reg(466) <= "10001111101111110000011110001000";
                        f_reg(467) <= "00010111110111111111111111111100";
                        f_reg(468) <= "00010000000000001111111100110110";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000001111100111";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
                  f_data <= f_data;
               end if;

            -- When attempting to write to memory
            elsif (i_write_enable = '1') then
               if (f_write = '0') then
                  f_write <= '1';
                  f_clk_count <= (others => '0');
                  f_timeout_flag <= '0';
                  case i_address is
                     when k_prog(1) =>
                        -- LUI R31 999
                        f_reg(1) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(2) =>
                        -- SRL R31 R31 16
                        f_reg(2) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(3) =>
                        -- LUI R1 -19413
                        f_reg(3) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(4) =>
                        -- SLTU R2 R1 R0
                        f_reg(4) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(5) =>
                        -- XORI R3 R2 -14645
                        f_reg(5) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(6) =>
                        -- SLLV R4 R2 R3
                        f_reg(6) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(7) =>
                        -- SLT R5 R1 R3
                        f_reg(7) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(8) =>
                        -- SLTIU R6 R4 29340
                        f_reg(8) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(9) =>
                        -- SLTIU R7 R6 -11769
                        f_reg(9) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(10) =>
                        -- XOR R8 R7 R7
                        f_reg(10) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(11) =>
                        -- ORI R9 R5 27837
                        f_reg(11) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(12) =>
                        -- SRLV R10 R5 R2
                        f_reg(12) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(13) =>
                        -- SLL R11 R7 18
                        f_reg(13) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(14) =>
                        -- SW R3 R0 1080
                        f_reg(14) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(15) =>
                        -- SUB R12 R2 R9
                        f_reg(15) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(16) =>
                        -- OR R13 R4 R0
                        f_reg(16) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(17) =>
                        -- ORI R14 R0 30369
                        f_reg(17) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(18) =>
                        -- SLT R15 R12 R13
                        f_reg(18) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(19) =>
                        -- SRLV R16 R15 R8
                        f_reg(19) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(20) =>
                        -- XOR R17 R2 R15
                        f_reg(20) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(21) =>
                        -- LUI R18 9669
                        f_reg(21) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(22) =>
                        -- SLL R19 R5 21
                        f_reg(22) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(23) =>
                        -- SLTU R20 R13 R14
                        f_reg(23) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(24) =>
                        -- SUBU R21 R2 R2
                        f_reg(24) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(25) =>
                        -- SLLV R14 R14 R3
                        f_reg(25) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(26) =>
                        -- ADDIU R22 R3 -26681
                        f_reg(26) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(27) =>
                        -- SRLV R23 R16 R22
                        f_reg(27) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(28) =>
                        -- ANDI R24 R20 32377
                        f_reg(28) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(29) =>
                        -- SUBU R25 R4 R24
                        f_reg(29) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(30) =>
                        -- SW R18 R0 1084
                        f_reg(30) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(31) =>
                        -- SRAV R26 R21 R9
                        f_reg(31) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(32) =>
                        -- ADDIU R27 R26 -11907
                        f_reg(32) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(33) =>
                        -- OR R28 R24 R10
                        f_reg(33) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(34) =>
                        -- ORI R29 R5 27080
                        f_reg(34) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(35) =>
                        -- SW R28 R0 1088
                        f_reg(35) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(36) =>
                        -- SRLV R30 R6 R23
                        f_reg(36) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(37) =>
                        -- OR R1 R26 R22
                        f_reg(37) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(38) =>
                        -- SW R28 R0 1092
                        f_reg(38) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(39) =>
                        -- ANDI R12 R30 -22366
                        f_reg(39) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(40) =>
                        -- SLT R8 R9 R29
                        f_reg(40) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(41) =>
                        -- XOR R4 R12 R4
                        f_reg(41) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(42) =>
                        -- SLT R15 R14 R27
                        f_reg(42) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(43) =>
                        -- SUBU R2 R11 R17
                        f_reg(43) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(44) =>
                        -- SRL R3 R12 5
                        f_reg(44) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(45) =>
                        -- SUB R16 R8 R19
                        f_reg(45) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(46) =>
                        -- XOR R20 R4 R7
                        f_reg(46) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(47) =>
                        -- ADDU R18 R2 R13
                        f_reg(47) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(48) =>
                        -- SLLV R21 R1 R7
                        f_reg(48) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(49) =>
                        -- SLTIU R10 R3 25015
                        f_reg(49) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(50) =>
                        -- NOR R5 R21 R25
                        f_reg(50) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(51) =>
                        -- NOP
                        f_reg(51) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(52) =>
                        -- SLTIU R6 R19 23581
                        f_reg(52) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(53) =>
                        -- SLLV R23 R5 R18
                        f_reg(53) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(54) =>
                        -- SLTI R26 R27 29940
                        f_reg(54) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(55) =>
                        -- SRL R22 R15 14
                        f_reg(55) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(56) =>
                        -- NOP
                        f_reg(56) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(57) =>
                        -- SW R19 R0 1096
                        f_reg(57) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(58) =>
                        -- ANDI R28 R26 -1792
                        f_reg(58) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(59) =>
                        -- NOR R9 R23 R20
                        f_reg(59) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(60) =>
                        -- LUI R29 -16537
                        f_reg(60) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(61) =>
                        -- SRAV R14 R16 R10
                        f_reg(61) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(62) =>
                        -- AND R11 R14 R6
                        f_reg(62) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(63) =>
                        -- NOP
                        f_reg(63) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(64) =>
                        -- SW R11 R0 1100
                        f_reg(64) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(65) =>
                        -- XOR R17 R22 R22
                        f_reg(65) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(66) =>
                        -- SW R30 R0 1104
                        f_reg(66) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(67) =>
                        -- SLL R12 R0 24
                        f_reg(67) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(68) =>
                        -- ADDIU R8 R29 8233
                        f_reg(68) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(69) =>
                        -- NOR R4 R17 R24
                        f_reg(69) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(70) =>
                        -- SRLV R2 R8 R13
                        f_reg(70) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(71) =>
                        -- NOP
                        f_reg(71) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(72) =>
                        -- XOR R1 R12 R28
                        f_reg(72) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(73) =>
                        -- SLLV R7 R1 R2
                        f_reg(73) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(74) =>
                        -- NOP
                        f_reg(74) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(75) =>
                        -- SW R9 R0 1108
                        f_reg(75) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(76) =>
                        -- SW R7 R0 1112
                        f_reg(76) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(77) =>
                        -- SW R4 R0 1116
                        f_reg(77) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(78) =>
                        -- ADDI R31 R31 -1
                        f_reg(78) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(79) =>
                        -- BGTZ R31 -76
                        f_reg(79) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(80) =>
                        -- BEQ R0 R0 454
                        f_reg(80) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(81) =>
                        -- LUI R30 999
                        f_reg(81) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(82) =>
                        -- LUI R31 999
                        f_reg(82) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(83) =>
                        -- SRL R30 R30 16
                        f_reg(83) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(84) =>
                        -- SRL R31 R31 16
                        f_reg(84) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(85) =>
                        -- LUI R1 -19413
                        f_reg(85) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(86) =>
                        -- LUI R15 -19413
                        f_reg(86) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(87) =>
                        -- SLTU R2 R1 R0
                        f_reg(87) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(88) =>
                        -- SLTU R16 R15 R0
                        f_reg(88) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(89) =>
                        -- XORI R3 R2 -14645
                        f_reg(89) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(90) =>
                        -- XORI R17 R16 -14645
                        f_reg(90) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(91) =>
                        -- SLLV R4 R2 R3
                        f_reg(91) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(92) =>
                        -- SLLV R18 R16 R17
                        f_reg(92) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(93) =>
                        -- SLT R5 R1 R3
                        f_reg(93) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(94) =>
                        -- SLT R19 R15 R17
                        f_reg(94) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(95) =>
                        -- SLTIU R6 R4 29340
                        f_reg(95) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(96) =>
                        -- SLTIU R20 R18 29340
                        f_reg(96) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(97) =>
                        -- SLTIU R7 R6 -11769
                        f_reg(97) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(98) =>
                        -- SLTIU R21 R20 -11769
                        f_reg(98) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(99) =>
                        -- XOR R8 R7 R7
                        f_reg(99) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(100) =>
                        -- XOR R22 R21 R21
                        f_reg(100) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(101) =>
                        -- ORI R9 R5 27837
                        f_reg(101) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(102) =>
                        -- ORI R23 R19 27837
                        f_reg(102) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(103) =>
                        -- SRLV R10 R5 R2
                        f_reg(103) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(104) =>
                        -- SRLV R24 R19 R16
                        f_reg(104) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(105) =>
                        -- SLL R11 R7 18
                        f_reg(105) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(106) =>
                        -- SLL R25 R21 18
                        f_reg(106) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(107) =>
                        -- BNE R3 R17 286
                        f_reg(107) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(108) =>
                        -- SW R3 R0 1080
                        f_reg(108) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(109) =>
                        -- SUB R12 R2 R9
                        f_reg(109) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(110) =>
                        -- SUB R26 R16 R23
                        f_reg(110) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(111) =>
                        -- OR R13 R4 R0
                        f_reg(111) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(112) =>
                        -- OR R27 R18 R0
                        f_reg(112) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(113) =>
                        -- ORI R14 R0 30369
                        f_reg(113) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(114) =>
                        -- ORI R28 R0 30369
                        f_reg(114) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(115) =>
                        -- SLT R1 R12 R13
                        f_reg(115) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(116) =>
                        -- SLT R15 R26 R27
                        f_reg(116) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(117) =>
                        -- SRLV R12 R1 R8
                        f_reg(117) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(118) =>
                        -- SRLV R26 R15 R22
                        f_reg(118) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(119) =>
                        -- XOR R8 R2 R1
                        f_reg(119) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(120) =>
                        -- XOR R22 R16 R15
                        f_reg(120) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(121) =>
                        -- LUI R1 9669
                        f_reg(121) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(122) =>
                        -- LUI R15 9669
                        f_reg(122) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(123) =>
                        -- BNE R13 R27 270
                        f_reg(123) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(124) =>
                        -- SW R13 R0 1120
                        f_reg(124) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(125) =>
                        -- SLL R13 R5 21
                        f_reg(125) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(126) =>
                        -- SLL R27 R19 21
                        f_reg(126) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(127) =>
                        -- BNE R13 R27 266
                        f_reg(127) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(128) =>
                        -- SW R13 R0 1124
                        f_reg(128) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(129) =>
                        -- LW R13 R0 1120
                        f_reg(129) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(130) =>
                        -- LW R27 R0 1120
                        f_reg(130) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(131) =>
                        -- BNE R13 R27 -2
                        f_reg(131) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(132) =>
                        -- BNE R7 R21 261
                        f_reg(132) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(133) =>
                        -- SW R7 R0 1128
                        f_reg(133) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(134) =>
                        -- SLTU R7 R13 R14
                        f_reg(134) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(135) =>
                        -- SLTU R21 R27 R28
                        f_reg(135) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(136) =>
                        -- BNE R13 R27 257
                        f_reg(136) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(137) =>
                        -- SW R13 R0 1132
                        f_reg(137) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(138) =>
                        -- SUBU R13 R2 R2
                        f_reg(138) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(139) =>
                        -- SUBU R27 R16 R16
                        f_reg(139) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(140) =>
                        -- SLLV R14 R14 R3
                        f_reg(140) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(141) =>
                        -- SLLV R28 R28 R17
                        f_reg(141) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(142) =>
                        -- ADDIU R2 R3 -26681
                        f_reg(142) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(143) =>
                        -- ADDIU R16 R17 -26681
                        f_reg(143) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(144) =>
                        -- SRLV R3 R12 R2
                        f_reg(144) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(145) =>
                        -- SRLV R17 R26 R16
                        f_reg(145) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(146) =>
                        -- ANDI R12 R7 32377
                        f_reg(146) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(147) =>
                        -- ANDI R26 R21 32377
                        f_reg(147) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(148) =>
                        -- SUBU R7 R4 R12
                        f_reg(148) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(149) =>
                        -- SUBU R21 R18 R26
                        f_reg(149) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(150) =>
                        -- BNE R1 R15 243
                        f_reg(150) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(151) =>
                        -- SW R1 R0 1084
                        f_reg(151) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(152) =>
                        -- SRAV R1 R13 R9
                        f_reg(152) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(153) =>
                        -- SRAV R15 R27 R23
                        f_reg(153) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(154) =>
                        -- ADDIU R13 R1 -11907
                        f_reg(154) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(155) =>
                        -- ADDIU R27 R15 -11907
                        f_reg(155) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(156) =>
                        -- BNE R13 R27 237
                        f_reg(156) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(157) =>
                        -- SW R13 R0 1136
                        f_reg(157) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(158) =>
                        -- OR R13 R12 R10
                        f_reg(158) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(159) =>
                        -- OR R27 R26 R24
                        f_reg(159) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(160) =>
                        -- ORI R10 R5 27080
                        f_reg(160) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(161) =>
                        -- ORI R24 R19 27080
                        f_reg(161) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(162) =>
                        -- BNE R13 R27 231
                        f_reg(162) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(163) =>
                        -- SW R13 R0 1088
                        f_reg(163) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(164) =>
                        -- SRLV R5 R6 R3
                        f_reg(164) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(165) =>
                        -- SRLV R19 R20 R17
                        f_reg(165) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(166) =>
                        -- OR R6 R1 R2
                        f_reg(166) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(167) =>
                        -- OR R20 R15 R16
                        f_reg(167) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(168) =>
                        -- BNE R13 R27 225
                        f_reg(168) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(169) =>
                        -- SW R13 R0 1092
                        f_reg(169) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(170) =>
                        -- ANDI R3 R5 -22366
                        f_reg(170) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(171) =>
                        -- ANDI R17 R19 -22366
                        f_reg(171) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(172) =>
                        -- SLT R1 R9 R10
                        f_reg(172) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(173) =>
                        -- SLT R15 R23 R24
                        f_reg(173) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(174) =>
                        -- XOR R4 R3 R4
                        f_reg(174) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(175) =>
                        -- XOR R18 R17 R18
                        f_reg(175) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(176) =>
                        -- LW R2 R0 1136
                        f_reg(176) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(177) =>
                        -- LW R16 R0 1136
                        f_reg(177) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(178) =>
                        -- BNE R2 R16 -2
                        f_reg(178) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(179) =>
                        -- SLT R13 R14 R2
                        f_reg(179) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(180) =>
                        -- SLT R27 R28 R16
                        f_reg(180) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(181) =>
                        -- SUBU R9 R11 R8
                        f_reg(181) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(182) =>
                        -- SUBU R23 R25 R22
                        f_reg(182) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(183) =>
                        -- SRL R10 R3 5
                        f_reg(183) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(184) =>
                        -- SRL R24 R17 5
                        f_reg(184) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(185) =>
                        -- LW R14 R0 1124
                        f_reg(185) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(186) =>
                        -- LW R28 R0 1124
                        f_reg(186) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(187) =>
                        -- BNE R14 R28 -2
                        f_reg(187) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(188) =>
                        -- SUB R11 R1 R14
                        f_reg(188) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(189) =>
                        -- SUB R25 R15 R28
                        f_reg(189) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(190) =>
                        -- LW R8 R0 1128
                        f_reg(190) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(191) =>
                        -- LW R22 R0 1128
                        f_reg(191) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(192) =>
                        -- BNE R8 R22 -2
                        f_reg(192) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(193) =>
                        -- XOR R3 R4 R8
                        f_reg(193) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(194) =>
                        -- XOR R17 R18 R22
                        f_reg(194) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(195) =>
                        -- LW R1 R0 1132
                        f_reg(195) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(196) =>
                        -- LW R15 R0 1132
                        f_reg(196) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(197) =>
                        -- BNE R1 R15 -2
                        f_reg(197) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(198) =>
                        -- ADDU R4 R9 R1
                        f_reg(198) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(199) =>
                        -- ADDU R18 R23 R15
                        f_reg(199) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(200) =>
                        -- SLLV R9 R6 R8
                        f_reg(200) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(201) =>
                        -- SLLV R23 R20 R22
                        f_reg(201) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(202) =>
                        -- SLTIU R6 R10 25015
                        f_reg(202) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(203) =>
                        -- SLTIU R20 R24 25015
                        f_reg(203) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(204) =>
                        -- NOR R8 R9 R7
                        f_reg(204) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(205) =>
                        -- NOR R22 R23 R21
                        f_reg(205) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(206) =>
                        -- NOP
                        f_reg(206) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(207) =>
                        -- NOP
                        f_reg(207) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(208) =>
                        -- SLTIU R10 R14 23581
                        f_reg(208) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(209) =>
                        -- SLTIU R24 R28 23581
                        f_reg(209) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(210) =>
                        -- SLLV R9 R8 R4
                        f_reg(210) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(211) =>
                        -- SLLV R23 R22 R18
                        f_reg(211) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(212) =>
                        -- SLTI R7 R2 29940
                        f_reg(212) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(213) =>
                        -- SLTI R21 R16 29940
                        f_reg(213) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(214) =>
                        -- SRL R8 R13 14
                        f_reg(214) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(215) =>
                        -- SRL R22 R27 14
                        f_reg(215) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(216) =>
                        -- NOP
                        f_reg(216) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(217) =>
                        -- NOP
                        f_reg(217) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(218) =>
                        -- BNE R14 R28 175
                        f_reg(218) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(219) =>
                        -- SW R14 R0 1096
                        f_reg(219) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(220) =>
                        -- ANDI R4 R7 -1792
                        f_reg(220) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(221) =>
                        -- ANDI R18 R21 -1792
                        f_reg(221) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(222) =>
                        -- NOR R2 R9 R3
                        f_reg(222) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(223) =>
                        -- NOR R16 R23 R17
                        f_reg(223) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(224) =>
                        -- LUI R13 -16537
                        f_reg(224) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(225) =>
                        -- LUI R27 -16537
                        f_reg(225) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(226) =>
                        -- SRAV R14 R11 R6
                        f_reg(226) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(227) =>
                        -- SRAV R28 R25 R20
                        f_reg(227) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(228) =>
                        -- AND R7 R14 R10
                        f_reg(228) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(229) =>
                        -- AND R21 R28 R24
                        f_reg(229) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(230) =>
                        -- NOP
                        f_reg(230) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(231) =>
                        -- NOP
                        f_reg(231) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(232) =>
                        -- BNE R7 R21 161
                        f_reg(232) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(233) =>
                        -- SW R7 R0 1100
                        f_reg(233) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(234) =>
                        -- XOR R9 R8 R8
                        f_reg(234) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(235) =>
                        -- XOR R23 R22 R22
                        f_reg(235) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(236) =>
                        -- BNE R5 R19 157
                        f_reg(236) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(237) =>
                        -- SW R5 R0 1104
                        f_reg(237) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(238) =>
                        -- SLL R3 R0 24
                        f_reg(238) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(239) =>
                        -- SLL R17 R0 24
                        f_reg(239) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(240) =>
                        -- ADDIU R11 R13 8233
                        f_reg(240) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(241) =>
                        -- ADDIU R25 R27 8233
                        f_reg(241) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(242) =>
                        -- NOR R6 R9 R12
                        f_reg(242) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(243) =>
                        -- NOR R20 R23 R26
                        f_reg(243) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(244) =>
                        -- SRLV R14 R11 R1
                        f_reg(244) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(245) =>
                        -- SRLV R28 R25 R15
                        f_reg(245) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(246) =>
                        -- NOP
                        f_reg(246) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(247) =>
                        -- NOP
                        f_reg(247) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(248) =>
                        -- XOR R10 R3 R4
                        f_reg(248) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(249) =>
                        -- XOR R24 R17 R18
                        f_reg(249) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(250) =>
                        -- SLLV R7 R10 R14
                        f_reg(250) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(251) =>
                        -- SLLV R21 R24 R28
                        f_reg(251) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(252) =>
                        -- NOP
                        f_reg(252) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(253) =>
                        -- NOP
                        f_reg(253) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(254) =>
                        -- BNE R2 R16 139
                        f_reg(254) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(255) =>
                        -- SW R2 R0 1108
                        f_reg(255) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(256) =>
                        -- BNE R7 R21 137
                        f_reg(256) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(257) =>
                        -- SW R7 R0 1112
                        f_reg(257) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(258) =>
                        -- BNE R6 R20 135
                        f_reg(258) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(259) =>
                        -- SW R6 R0 1116
                        f_reg(259) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(260) =>
                        -- ADDI R29 R30 -250
                        f_reg(260) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(261) =>
                        -- BEQ R29 R0 25
                        f_reg(261) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(262) =>
                        -- ADDI R29 R30 -500
                        f_reg(262) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(263) =>
                        -- BEQ R29 R0 23
                        f_reg(263) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(264) =>
                        -- ADDI R29 R30 -750
                        f_reg(264) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(265) =>
                        -- BEQ R29 R0 21
                        f_reg(265) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(266) =>
                        -- ADDI R30 R30 -1
                        f_reg(266) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(267) =>
                        -- ADDI R31 R31 -1
                        f_reg(267) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(268) =>
                        -- BNE R30 R31 125
                        f_reg(268) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(269) =>
                        -- BGTZ R31 -184
                        f_reg(269) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(270) =>
                        -- BEQ R0 R0 264
                        f_reg(270) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(271) =>
                        -- NOP
                        f_reg(271) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(272) =>
                        -- NOP
                        f_reg(272) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(273) =>
                        -- NOP
                        f_reg(273) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(274) =>
                        -- NOP
                        f_reg(274) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(275) =>
                        -- NOP
                        f_reg(275) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(276) =>
                        -- NOP
                        f_reg(276) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(277) =>
                        -- NOP
                        f_reg(277) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(278) =>
                        -- NOP
                        f_reg(278) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(279) =>
                        -- NOP
                        f_reg(279) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(280) =>
                        -- NOP
                        f_reg(280) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(281) =>
                        -- NOP
                        f_reg(281) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(282) =>
                        -- NOP
                        f_reg(282) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(283) =>
                        -- NOP
                        f_reg(283) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(284) =>
                        -- NOP
                        f_reg(284) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(285) =>
                        -- NOP
                        f_reg(285) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(286) =>
                        -- LW R29 R0 1992
                        f_reg(286) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(287) =>
                        -- BGTZ R29 3
                        f_reg(287) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(288) =>
                        -- ADDI R29 R0 60
                        f_reg(288) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(289) =>
                        -- BEQ R0 R0 2
                        f_reg(289) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(290) =>
                        -- ADDI R29 R0 0
                        f_reg(290) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(291) =>
                        -- BNE R1 R15 102
                        f_reg(291) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(292) =>
                        -- SW R1 R29 1872
                        f_reg(292) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(293) =>
                        -- LW R29 R0 1992
                        f_reg(293) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(294) =>
                        -- BGTZ R29 3
                        f_reg(294) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(295) =>
                        -- ADDI R29 R0 60
                        f_reg(295) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(296) =>
                        -- BEQ R0 R0 2
                        f_reg(296) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(297) =>
                        -- ADDI R29 R0 0
                        f_reg(297) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(298) =>
                        -- BNE R2 R16 95
                        f_reg(298) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(299) =>
                        -- SW R2 R29 1876
                        f_reg(299) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(300) =>
                        -- LW R29 R0 1992
                        f_reg(300) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(301) =>
                        -- BGTZ R29 3
                        f_reg(301) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(302) =>
                        -- ADDI R29 R0 60
                        f_reg(302) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(303) =>
                        -- BEQ R0 R0 2
                        f_reg(303) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(304) =>
                        -- ADDI R29 R0 0
                        f_reg(304) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(305) =>
                        -- BNE R3 R17 88
                        f_reg(305) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(306) =>
                        -- SW R3 R29 1880
                        f_reg(306) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(307) =>
                        -- LW R29 R0 1992
                        f_reg(307) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(308) =>
                        -- BGTZ R29 3
                        f_reg(308) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(309) =>
                        -- ADDI R29 R0 60
                        f_reg(309) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(310) =>
                        -- BEQ R0 R0 2
                        f_reg(310) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(311) =>
                        -- ADDI R29 R0 0
                        f_reg(311) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(312) =>
                        -- BNE R4 R18 81
                        f_reg(312) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(313) =>
                        -- SW R4 R29 1884
                        f_reg(313) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(314) =>
                        -- LW R29 R0 1992
                        f_reg(314) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(315) =>
                        -- BGTZ R29 3
                        f_reg(315) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(316) =>
                        -- ADDI R29 R0 60
                        f_reg(316) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(317) =>
                        -- BEQ R0 R0 2
                        f_reg(317) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(318) =>
                        -- ADDI R29 R0 0
                        f_reg(318) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(319) =>
                        -- BNE R5 R19 74
                        f_reg(319) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(320) =>
                        -- SW R5 R29 1888
                        f_reg(320) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(321) =>
                        -- LW R29 R0 1992
                        f_reg(321) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(322) =>
                        -- BGTZ R29 3
                        f_reg(322) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(323) =>
                        -- ADDI R29 R0 60
                        f_reg(323) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(324) =>
                        -- BEQ R0 R0 2
                        f_reg(324) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(325) =>
                        -- ADDI R29 R0 0
                        f_reg(325) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(326) =>
                        -- BNE R6 R20 67
                        f_reg(326) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(327) =>
                        -- SW R6 R29 1892
                        f_reg(327) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(328) =>
                        -- LW R29 R0 1992
                        f_reg(328) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(329) =>
                        -- BGTZ R29 3
                        f_reg(329) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(330) =>
                        -- ADDI R29 R0 60
                        f_reg(330) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(331) =>
                        -- BEQ R0 R0 2
                        f_reg(331) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(332) =>
                        -- ADDI R29 R0 0
                        f_reg(332) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(333) =>
                        -- BNE R7 R21 60
                        f_reg(333) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(334) =>
                        -- SW R7 R29 1896
                        f_reg(334) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(335) =>
                        -- LW R29 R0 1992
                        f_reg(335) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(336) =>
                        -- BGTZ R29 3
                        f_reg(336) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(337) =>
                        -- ADDI R29 R0 60
                        f_reg(337) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(338) =>
                        -- BEQ R0 R0 2
                        f_reg(338) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(339) =>
                        -- ADDI R29 R0 0
                        f_reg(339) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(340) =>
                        -- BNE R8 R22 53
                        f_reg(340) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(341) =>
                        -- SW R8 R29 1900
                        f_reg(341) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(342) =>
                        -- LW R29 R0 1992
                        f_reg(342) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(343) =>
                        -- BGTZ R29 3
                        f_reg(343) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(344) =>
                        -- ADDI R29 R0 60
                        f_reg(344) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(345) =>
                        -- BEQ R0 R0 2
                        f_reg(345) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(346) =>
                        -- ADDI R29 R0 0
                        f_reg(346) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(347) =>
                        -- BNE R9 R23 46
                        f_reg(347) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(348) =>
                        -- SW R9 R29 1904
                        f_reg(348) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(349) =>
                        -- LW R29 R0 1992
                        f_reg(349) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(350) =>
                        -- BGTZ R29 3
                        f_reg(350) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(351) =>
                        -- ADDI R29 R0 60
                        f_reg(351) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(352) =>
                        -- BEQ R0 R0 2
                        f_reg(352) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(353) =>
                        -- ADDI R29 R0 0
                        f_reg(353) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(354) =>
                        -- BNE R10 R24 39
                        f_reg(354) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(355) =>
                        -- SW R10 R29 1908
                        f_reg(355) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(356) =>
                        -- LW R29 R0 1992
                        f_reg(356) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(357) =>
                        -- BGTZ R29 3
                        f_reg(357) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(358) =>
                        -- ADDI R29 R0 60
                        f_reg(358) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(359) =>
                        -- BEQ R0 R0 2
                        f_reg(359) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(360) =>
                        -- ADDI R29 R0 0
                        f_reg(360) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(361) =>
                        -- BNE R11 R25 32
                        f_reg(361) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(362) =>
                        -- SW R11 R29 1912
                        f_reg(362) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(363) =>
                        -- LW R29 R0 1992
                        f_reg(363) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(364) =>
                        -- BGTZ R29 3
                        f_reg(364) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(365) =>
                        -- ADDI R29 R0 60
                        f_reg(365) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(366) =>
                        -- BEQ R0 R0 2
                        f_reg(366) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(367) =>
                        -- ADDI R29 R0 0
                        f_reg(367) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(368) =>
                        -- BNE R12 R26 25
                        f_reg(368) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(369) =>
                        -- SW R12 R29 1916
                        f_reg(369) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(370) =>
                        -- LW R29 R0 1992
                        f_reg(370) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(371) =>
                        -- BGTZ R29 3
                        f_reg(371) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(372) =>
                        -- ADDI R29 R0 60
                        f_reg(372) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(373) =>
                        -- BEQ R0 R0 2
                        f_reg(373) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(374) =>
                        -- ADDI R29 R0 0
                        f_reg(374) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(375) =>
                        -- BNE R13 R27 18
                        f_reg(375) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(376) =>
                        -- SW R13 R29 1920
                        f_reg(376) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(377) =>
                        -- LW R29 R0 1992
                        f_reg(377) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(378) =>
                        -- BGTZ R29 3
                        f_reg(378) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(379) =>
                        -- ADDI R29 R0 60
                        f_reg(379) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(380) =>
                        -- BEQ R0 R0 2
                        f_reg(380) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(381) =>
                        -- ADDI R29 R0 0
                        f_reg(381) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(382) =>
                        -- BNE R14 R28 11
                        f_reg(382) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(383) =>
                        -- SW R14 R29 1924
                        f_reg(383) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(384) =>
                        -- LW R29 R0 1992
                        f_reg(384) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(385) =>
                        -- BGTZ R29 3
                        f_reg(385) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(386) =>
                        -- ADDI R29 R0 60
                        f_reg(386) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(387) =>
                        -- BEQ R0 R0 2
                        f_reg(387) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(388) =>
                        -- ADDI R29 R0 0
                        f_reg(388) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(389) =>
                        -- BNE R30 R31 4
                        f_reg(389) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(390) =>
                        -- SW R30 R29 1928
                        f_reg(390) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(391) =>
                        -- SW R29 R0 1992
                        f_reg(391) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(392) =>
                        -- BEQ R0 R0 -126
                        f_reg(392) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(393) =>
                        -- LW R29 R0 1992
                        f_reg(393) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(394) =>
                        -- LW R1 R29 1872
                        f_reg(394) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(395) =>
                        -- LW R29 R0 1992
                        f_reg(395) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(396) =>
                        -- LW R15 R29 1872
                        f_reg(396) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(397) =>
                        -- BNE R1 R15 -4
                        f_reg(397) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(398) =>
                        -- LW R29 R0 1992
                        f_reg(398) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(399) =>
                        -- LW R2 R29 1876
                        f_reg(399) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(400) =>
                        -- LW R29 R0 1992
                        f_reg(400) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(401) =>
                        -- LW R16 R29 1876
                        f_reg(401) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(402) =>
                        -- BNE R2 R16 -4
                        f_reg(402) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(403) =>
                        -- LW R29 R0 1992
                        f_reg(403) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(404) =>
                        -- LW R3 R29 1880
                        f_reg(404) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(405) =>
                        -- LW R29 R0 1992
                        f_reg(405) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(406) =>
                        -- LW R17 R29 1880
                        f_reg(406) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(407) =>
                        -- BNE R3 R17 -4
                        f_reg(407) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(408) =>
                        -- LW R29 R0 1992
                        f_reg(408) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(409) =>
                        -- LW R4 R29 1884
                        f_reg(409) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(410) =>
                        -- LW R29 R0 1992
                        f_reg(410) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(411) =>
                        -- LW R18 R29 1884
                        f_reg(411) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(412) =>
                        -- BNE R4 R18 -4
                        f_reg(412) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(413) =>
                        -- LW R29 R0 1992
                        f_reg(413) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(414) =>
                        -- LW R5 R29 1888
                        f_reg(414) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(415) =>
                        -- LW R29 R0 1992
                        f_reg(415) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(416) =>
                        -- LW R19 R29 1888
                        f_reg(416) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(417) =>
                        -- BNE R5 R19 -4
                        f_reg(417) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(418) =>
                        -- LW R29 R0 1992
                        f_reg(418) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(419) =>
                        -- LW R6 R29 1892
                        f_reg(419) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(420) =>
                        -- LW R29 R0 1992
                        f_reg(420) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(421) =>
                        -- LW R20 R29 1892
                        f_reg(421) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(422) =>
                        -- BNE R6 R20 -4
                        f_reg(422) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(423) =>
                        -- LW R29 R0 1992
                        f_reg(423) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(424) =>
                        -- LW R7 R29 1896
                        f_reg(424) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(425) =>
                        -- LW R29 R0 1992
                        f_reg(425) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(426) =>
                        -- LW R21 R29 1896
                        f_reg(426) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(427) =>
                        -- BNE R7 R21 -4
                        f_reg(427) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(428) =>
                        -- LW R29 R0 1992
                        f_reg(428) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(429) =>
                        -- LW R8 R29 1900
                        f_reg(429) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(430) =>
                        -- LW R29 R0 1992
                        f_reg(430) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(431) =>
                        -- LW R22 R29 1900
                        f_reg(431) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(432) =>
                        -- BNE R8 R22 -4
                        f_reg(432) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(433) =>
                        -- LW R29 R0 1992
                        f_reg(433) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(434) =>
                        -- LW R9 R29 1904
                        f_reg(434) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(435) =>
                        -- LW R29 R0 1992
                        f_reg(435) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(436) =>
                        -- LW R23 R29 1904
                        f_reg(436) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(437) =>
                        -- BNE R9 R23 -4
                        f_reg(437) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(438) =>
                        -- LW R29 R0 1992
                        f_reg(438) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(439) =>
                        -- LW R10 R29 1908
                        f_reg(439) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(440) =>
                        -- LW R29 R0 1992
                        f_reg(440) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(441) =>
                        -- LW R24 R29 1908
                        f_reg(441) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(442) =>
                        -- BNE R10 R24 -4
                        f_reg(442) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(443) =>
                        -- LW R29 R0 1992
                        f_reg(443) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(444) =>
                        -- LW R11 R29 1912
                        f_reg(444) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(445) =>
                        -- LW R29 R0 1992
                        f_reg(445) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(446) =>
                        -- LW R25 R29 1912
                        f_reg(446) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(447) =>
                        -- BNE R11 R25 -4
                        f_reg(447) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(448) =>
                        -- LW R29 R0 1992
                        f_reg(448) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(449) =>
                        -- LW R12 R29 1916
                        f_reg(449) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(450) =>
                        -- LW R29 R0 1992
                        f_reg(450) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(451) =>
                        -- LW R26 R29 1916
                        f_reg(451) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(452) =>
                        -- BNE R12 R26 -4
                        f_reg(452) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(453) =>
                        -- LW R29 R0 1992
                        f_reg(453) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(454) =>
                        -- LW R13 R29 1920
                        f_reg(454) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(455) =>
                        -- LW R29 R0 1992
                        f_reg(455) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(456) =>
                        -- LW R27 R29 1920
                        f_reg(456) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(457) =>
                        -- BNE R13 R27 -4
                        f_reg(457) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(458) =>
                        -- LW R29 R0 1992
                        f_reg(458) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(459) =>
                        -- LW R14 R29 1924
                        f_reg(459) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(460) =>
                        -- LW R29 R0 1992
                        f_reg(460) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(461) =>
                        -- LW R28 R29 1924
                        f_reg(461) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(462) =>
                        -- BNE R14 R28 -4
                        f_reg(462) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(463) =>
                        -- LW R29 R0 1992
                        f_reg(463) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(464) =>
                        -- LW R30 R29 1928
                        f_reg(464) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(465) =>
                        -- LW R29 R0 1992
                        f_reg(465) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(466) =>
                        -- LW R31 R29 1928
                        f_reg(466) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(467) =>
                        -- BNE R30 R31 -4
                        f_reg(467) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(468) =>
                        -- BEQ R0 R0 -202
                        f_reg(468) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(469) =>
                        -- NOP
                        f_reg(469) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(470) =>
                        -- NOP
                        f_reg(470) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(471) =>
                        -- NOP
                        f_reg(471) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(472) =>
                        -- NOP
                        f_reg(472) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(473) =>
                        -- NOP
                        f_reg(473) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(474) =>
                        -- NOP
                        f_reg(474) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(475) =>
                        -- NOP
                        f_reg(475) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(476) =>
                        -- NOP
                        f_reg(476) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(477) =>
                        -- NOP
                        f_reg(477) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(478) =>
                        -- NOP
                        f_reg(478) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(479) =>
                        -- NOP
                        f_reg(479) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(480) =>
                        -- NOP
                        f_reg(480) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(481) =>
                        -- NOP
                        f_reg(481) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(482) =>
                        -- NOP
                        f_reg(482) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(483) =>
                        -- NOP
                        f_reg(483) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(484) =>
                        -- NOP
                        f_reg(484) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(485) =>
                        -- NOP
                        f_reg(485) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(486) =>
                        -- NOP
                        f_reg(486) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(487) =>
                        -- NOP
                        f_reg(487) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(488) =>
                        -- NOP
                        f_reg(488) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(489) =>
                        -- NOP
                        f_reg(489) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(490) =>
                        -- NOP
                        f_reg(490) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(491) =>
                        -- NOP
                        f_reg(491) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(492) =>
                        -- NOP
                        f_reg(492) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(493) =>
                        -- NOP
                        f_reg(493) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(494) =>
                        -- NOP
                        f_reg(494) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(495) =>
                        -- NOP
                        f_reg(495) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(496) =>
                        -- NOP
                        f_reg(496) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(497) =>
                        -- NOP
                        f_reg(497) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(498) =>
                        -- NOP
                        f_reg(498) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(499) =>
                        -- NOP
                        f_reg(499) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(500) =>
                        -- NOP
                        f_reg(500) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(501) =>
                        -- NOP
                        f_reg(501) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(502) =>
                        -- NOP
                        f_reg(502) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(503) =>
                        -- NOP
                        f_reg(503) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(504) =>
                        -- NOP
                        f_reg(504) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(505) =>
                        -- NOP
                        f_reg(505) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(506) =>
                        -- NOP
                        f_reg(506) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(507) =>
                        -- NOP
                        f_reg(507) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(508) =>
                        -- NOP
                        f_reg(508) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(509) =>
                        -- NOP
                        f_reg(509) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(510) =>
                        -- NOP
                        f_reg(510) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(511) =>
                        -- NOP
                        f_reg(511) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(512) =>
                        -- NOP
                        f_reg(512) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(513) =>
                        -- NOP
                        f_reg(513) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(514) =>
                        -- NOP
                        f_reg(514) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(515) =>
                        -- NOP
                        f_reg(515) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(516) =>
                        -- NOP
                        f_reg(516) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(517) =>
                        -- NOP
                        f_reg(517) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(518) =>
                        -- NOP
                        f_reg(518) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(519) =>
                        -- NOP
                        f_reg(519) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(520) =>
                        -- NOP
                        f_reg(520) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(521) =>
                        -- NOP
                        f_reg(521) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(522) =>
                        -- NOP
                        f_reg(522) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(523) =>
                        -- NOP
                        f_reg(523) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(524) =>
                        -- NOP
                        f_reg(524) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(525) =>
                        -- NOP
                        f_reg(525) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(526) =>
                        -- NOP
                        f_reg(526) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(527) =>
                        -- NOP
                        f_reg(527) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(528) =>
                        -- NOP
                        f_reg(528) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(529) =>
                        -- NOP
                        f_reg(529) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(530) =>
                        -- NOP
                        f_reg(530) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(531) =>
                        -- NOP
                        f_reg(531) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(532) =>
                        -- NOP
                        f_reg(532) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(533) =>
                        -- NOP
                        f_reg(533) <= i_data;
                        f_MEM_READY <= '1';
                     when k_prog(534) =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011011010000101011";
                        f_reg(4) <= "00000000001000000001000000101011";
                        f_reg(5) <= "00111000010000111100011011001011";
                        f_reg(6) <= "00000000011000100010000000000100";
                        f_reg(7) <= "00000000001000110010100000101010";
                        f_reg(8) <= "00101100100001100111001010011100";
                        f_reg(9) <= "00101100110001111101001000000111";
                        f_reg(10) <= "00000000111001110100000000100110";
                        f_reg(11) <= "00110100101010010110110010111101";
                        f_reg(12) <= "00000000010001010101000000000110";
                        f_reg(13) <= "00000000000001110101110010000000";
                        f_reg(14) <= "10101100000000110000010000111000";
                        f_reg(15) <= "00000000010010010110000000100010";
                        f_reg(16) <= "00000000100000000110100000100101";
                        f_reg(17) <= "00110100000011100111011010100001";
                        f_reg(18) <= "00000001100011010111100000101010";
                        f_reg(19) <= "00000001000011111000000000000110";
                        f_reg(20) <= "00000000010011111000100000100110";
                        f_reg(21) <= "00111100000100100010010111000101";
                        f_reg(22) <= "00000000000001011001110101000000";
                        f_reg(23) <= "00000001101011101010000000101011";
                        f_reg(24) <= "00000000010000101010100000100011";
                        f_reg(25) <= "00000000011011100111000000000100";
                        f_reg(26) <= "00100100011101101001011111000111";
                        f_reg(27) <= "00000010110100001011100000000110";
                        f_reg(28) <= "00110010100110000111111001111001";
                        f_reg(29) <= "00000000100110001100100000100011";
                        f_reg(30) <= "10101100000100100000010000111100";
                        f_reg(31) <= "00000001001101011101000000000111";
                        f_reg(32) <= "00100111010110111101000101111101";
                        f_reg(33) <= "00000011000010101110000000100101";
                        f_reg(34) <= "00110100101111010110100111001000";
                        f_reg(35) <= "10101100000111000000010001000000";
                        f_reg(36) <= "00000010111001101111000000000110";
                        f_reg(37) <= "00000011010101100000100000100101";
                        f_reg(38) <= "10101100000111000000010001000100";
                        f_reg(39) <= "00110011110011001010100010100010";
                        f_reg(40) <= "00000001001111010100000000101010";
                        f_reg(41) <= "00000001100001000010000000100110";
                        f_reg(42) <= "00000001110110110111100000101010";
                        f_reg(43) <= "00000001011100010001000000100011";
                        f_reg(44) <= "00000000000011000001100101000010";
                        f_reg(45) <= "00000001000100111000000000100010";
                        f_reg(46) <= "00000000100001111010000000100110";
                        f_reg(47) <= "00000000010011011001000000100001";
                        f_reg(48) <= "00000000111000011010100000000100";
                        f_reg(49) <= "00101100011010100110000110110111";
                        f_reg(50) <= "00000010101110010010100000100111";
                        f_reg(51) <= "00000000000000000000000000000000";
                        f_reg(52) <= "00101110011001100101110000011101";
                        f_reg(53) <= "00000010010001011011100000000100";
                        f_reg(54) <= "00101011011110100111010011110100";
                        f_reg(55) <= "00000000000011111011001110000010";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "10101100000100110000010001001000";
                        f_reg(58) <= "00110011010111001111100100000000";
                        f_reg(59) <= "00000010111101000100100000100111";
                        f_reg(60) <= "00111100000111011011111101100111";
                        f_reg(61) <= "00000001010100000111000000000111";
                        f_reg(62) <= "00000001110001100101100000100100";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000010110000010001001100";
                        f_reg(65) <= "00000010110101101000100000100110";
                        f_reg(66) <= "10101100000111100000010001010000";
                        f_reg(67) <= "00000000000000000110011000000000";
                        f_reg(68) <= "00100111101010000010000000101001";
                        f_reg(69) <= "00000010001110000010000000100111";
                        f_reg(70) <= "00000001101010000001000000000110";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000001100111000000100000100110";
                        f_reg(73) <= "00000000010000010011100000000100";
                        f_reg(74) <= "00000000000000000000000000000000";
                        f_reg(75) <= "10101100000010010000010001010100";
                        f_reg(76) <= "10101100000001110000010001011000";
                        f_reg(77) <= "10101100000001000000010001011100";
                        f_reg(78) <= "00100011111111111111111111111111";
                        f_reg(79) <= "00011111111000001111111110110100";
                        f_reg(80) <= "00010000000000000000000111000110";
                        f_reg(81) <= "00111100000111100000001111100111";
                        f_reg(82) <= "00111100000111110000001111100111";
                        f_reg(83) <= "00000000000111101111010000000010";
                        f_reg(84) <= "00000000000111111111110000000010";
                        f_reg(85) <= "00111100000000011011010000101011";
                        f_reg(86) <= "00111100000011111011010000101011";
                        f_reg(87) <= "00000000001000000001000000101011";
                        f_reg(88) <= "00000001111000001000000000101011";
                        f_reg(89) <= "00111000010000111100011011001011";
                        f_reg(90) <= "00111010000100011100011011001011";
                        f_reg(91) <= "00000000011000100010000000000100";
                        f_reg(92) <= "00000010001100001001000000000100";
                        f_reg(93) <= "00000000001000110010100000101010";
                        f_reg(94) <= "00000001111100011001100000101010";
                        f_reg(95) <= "00101100100001100111001010011100";
                        f_reg(96) <= "00101110010101000111001010011100";
                        f_reg(97) <= "00101100110001111101001000000111";
                        f_reg(98) <= "00101110100101011101001000000111";
                        f_reg(99) <= "00000000111001110100000000100110";
                        f_reg(100) <= "00000010101101011011000000100110";
                        f_reg(101) <= "00110100101010010110110010111101";
                        f_reg(102) <= "00110110011101110110110010111101";
                        f_reg(103) <= "00000000010001010101000000000110";
                        f_reg(104) <= "00000010000100111100000000000110";
                        f_reg(105) <= "00000000000001110101110010000000";
                        f_reg(106) <= "00000000000101011100110010000000";
                        f_reg(107) <= "00010100011100010000000100011110";
                        f_reg(108) <= "10101100000000110000010000111000";
                        f_reg(109) <= "00000000010010010110000000100010";
                        f_reg(110) <= "00000010000101111101000000100010";
                        f_reg(111) <= "00000000100000000110100000100101";
                        f_reg(112) <= "00000010010000001101100000100101";
                        f_reg(113) <= "00110100000011100111011010100001";
                        f_reg(114) <= "00110100000111000111011010100001";
                        f_reg(115) <= "00000001100011010000100000101010";
                        f_reg(116) <= "00000011010110110111100000101010";
                        f_reg(117) <= "00000001000000010110000000000110";
                        f_reg(118) <= "00000010110011111101000000000110";
                        f_reg(119) <= "00000000010000010100000000100110";
                        f_reg(120) <= "00000010000011111011000000100110";
                        f_reg(121) <= "00111100000000010010010111000101";
                        f_reg(122) <= "00111100000011110010010111000101";
                        f_reg(123) <= "00010101101110110000000100001110";
                        f_reg(124) <= "10101100000011010000010001100000";
                        f_reg(125) <= "00000000000001010110110101000000";
                        f_reg(126) <= "00000000000100111101110101000000";
                        f_reg(127) <= "00010101101110110000000100001010";
                        f_reg(128) <= "10101100000011010000010001100100";
                        f_reg(129) <= "10001100000011010000010001100000";
                        f_reg(130) <= "10001100000110110000010001100000";
                        f_reg(131) <= "00010101101110111111111111111110";
                        f_reg(132) <= "00010100111101010000000100000101";
                        f_reg(133) <= "10101100000001110000010001101000";
                        f_reg(134) <= "00000001101011100011100000101011";
                        f_reg(135) <= "00000011011111001010100000101011";
                        f_reg(136) <= "00010101101110110000000100000001";
                        f_reg(137) <= "10101100000011010000010001101100";
                        f_reg(138) <= "00000000010000100110100000100011";
                        f_reg(139) <= "00000010000100001101100000100011";
                        f_reg(140) <= "00000000011011100111000000000100";
                        f_reg(141) <= "00000010001111001110000000000100";
                        f_reg(142) <= "00100100011000101001011111000111";
                        f_reg(143) <= "00100110001100001001011111000111";
                        f_reg(144) <= "00000000010011000001100000000110";
                        f_reg(145) <= "00000010000110101000100000000110";
                        f_reg(146) <= "00110000111011000111111001111001";
                        f_reg(147) <= "00110010101110100111111001111001";
                        f_reg(148) <= "00000000100011000011100000100011";
                        f_reg(149) <= "00000010010110101010100000100011";
                        f_reg(150) <= "00010100001011110000000011110011";
                        f_reg(151) <= "10101100000000010000010000111100";
                        f_reg(152) <= "00000001001011010000100000000111";
                        f_reg(153) <= "00000010111110110111100000000111";
                        f_reg(154) <= "00100100001011011101000101111101";
                        f_reg(155) <= "00100101111110111101000101111101";
                        f_reg(156) <= "00010101101110110000000011101101";
                        f_reg(157) <= "10101100000011010000010001110000";
                        f_reg(158) <= "00000001100010100110100000100101";
                        f_reg(159) <= "00000011010110001101100000100101";
                        f_reg(160) <= "00110100101010100110100111001000";
                        f_reg(161) <= "00110110011110000110100111001000";
                        f_reg(162) <= "00010101101110110000000011100111";
                        f_reg(163) <= "10101100000011010000010001000000";
                        f_reg(164) <= "00000000011001100010100000000110";
                        f_reg(165) <= "00000010001101001001100000000110";
                        f_reg(166) <= "00000000001000100011000000100101";
                        f_reg(167) <= "00000001111100001010000000100101";
                        f_reg(168) <= "00010101101110110000000011100001";
                        f_reg(169) <= "10101100000011010000010001000100";
                        f_reg(170) <= "00110000101000111010100010100010";
                        f_reg(171) <= "00110010011100011010100010100010";
                        f_reg(172) <= "00000001001010100000100000101010";
                        f_reg(173) <= "00000010111110000111100000101010";
                        f_reg(174) <= "00000000011001000010000000100110";
                        f_reg(175) <= "00000010001100101001000000100110";
                        f_reg(176) <= "10001100000000100000010001110000";
                        f_reg(177) <= "10001100000100000000010001110000";
                        f_reg(178) <= "00010100010100001111111111111110";
                        f_reg(179) <= "00000001110000100110100000101010";
                        f_reg(180) <= "00000011100100001101100000101010";
                        f_reg(181) <= "00000001011010000100100000100011";
                        f_reg(182) <= "00000011001101101011100000100011";
                        f_reg(183) <= "00000000000000110101000101000010";
                        f_reg(184) <= "00000000000100011100000101000010";
                        f_reg(185) <= "10001100000011100000010001100100";
                        f_reg(186) <= "10001100000111000000010001100100";
                        f_reg(187) <= "00010101110111001111111111111110";
                        f_reg(188) <= "00000000001011100101100000100010";
                        f_reg(189) <= "00000001111111001100100000100010";
                        f_reg(190) <= "10001100000010000000010001101000";
                        f_reg(191) <= "10001100000101100000010001101000";
                        f_reg(192) <= "00010101000101101111111111111110";
                        f_reg(193) <= "00000000100010000001100000100110";
                        f_reg(194) <= "00000010010101101000100000100110";
                        f_reg(195) <= "10001100000000010000010001101100";
                        f_reg(196) <= "10001100000011110000010001101100";
                        f_reg(197) <= "00010100001011111111111111111110";
                        f_reg(198) <= "00000001001000010010000000100001";
                        f_reg(199) <= "00000010111011111001000000100001";
                        f_reg(200) <= "00000001000001100100100000000100";
                        f_reg(201) <= "00000010110101001011100000000100";
                        f_reg(202) <= "00101101010001100110000110110111";
                        f_reg(203) <= "00101111000101000110000110110111";
                        f_reg(204) <= "00000001001001110100000000100111";
                        f_reg(205) <= "00000010111101011011000000100111";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101101110010100101110000011101";
                        f_reg(209) <= "00101111100110000101110000011101";
                        f_reg(210) <= "00000000100010000100100000000100";
                        f_reg(211) <= "00000010010101101011100000000100";
                        f_reg(212) <= "00101000010001110111010011110100";
                        f_reg(213) <= "00101010000101010111010011110100";
                        f_reg(214) <= "00000000000011010100001110000010";
                        f_reg(215) <= "00000000000110111011001110000010";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "00010101110111000000000010101111";
                        f_reg(219) <= "10101100000011100000010001001000";
                        f_reg(220) <= "00110000111001001111100100000000";
                        f_reg(221) <= "00110010101100101111100100000000";
                        f_reg(222) <= "00000001001000110001000000100111";
                        f_reg(223) <= "00000010111100011000000000100111";
                        f_reg(224) <= "00111100000011011011111101100111";
                        f_reg(225) <= "00111100000110111011111101100111";
                        f_reg(226) <= "00000000110010110111000000000111";
                        f_reg(227) <= "00000010100110011110000000000111";
                        f_reg(228) <= "00000001110010100011100000100100";
                        f_reg(229) <= "00000011100110001010100000100100";
                        f_reg(230) <= "00000000000000000000000000000000";
                        f_reg(231) <= "00000000000000000000000000000000";
                        f_reg(232) <= "00010100111101010000000010100001";
                        f_reg(233) <= "10101100000001110000010001001100";
                        f_reg(234) <= "00000001000010000100100000100110";
                        f_reg(235) <= "00000010110101101011100000100110";
                        f_reg(236) <= "00010100101100110000000010011101";
                        f_reg(237) <= "10101100000001010000010001010000";
                        f_reg(238) <= "00000000000000000001111000000000";
                        f_reg(239) <= "00000000000000001000111000000000";
                        f_reg(240) <= "00100101101010110010000000101001";
                        f_reg(241) <= "00100111011110010010000000101001";
                        f_reg(242) <= "00000001001011000011000000100111";
                        f_reg(243) <= "00000010111110101010000000100111";
                        f_reg(244) <= "00000000001010110111000000000110";
                        f_reg(245) <= "00000001111110011110000000000110";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00000000011001000101000000100110";
                        f_reg(249) <= "00000010001100101100000000100110";
                        f_reg(250) <= "00000001110010100011100000000100";
                        f_reg(251) <= "00000011100110001010100000000100";
                        f_reg(252) <= "00000000000000000000000000000000";
                        f_reg(253) <= "00000000000000000000000000000000";
                        f_reg(254) <= "00010100010100000000000010001011";
                        f_reg(255) <= "10101100000000100000010001010100";
                        f_reg(256) <= "00010100111101010000000010001001";
                        f_reg(257) <= "10101100000001110000010001011000";
                        f_reg(258) <= "00010100110101000000000010000111";
                        f_reg(259) <= "10101100000001100000010001011100";
                        f_reg(260) <= "00100011110111011111111100000110";
                        f_reg(261) <= "00010011101000000000000000011001";
                        f_reg(262) <= "00100011110111011111111000001100";
                        f_reg(263) <= "00010011101000000000000000010111";
                        f_reg(264) <= "00100011110111011111110100010010";
                        f_reg(265) <= "00010011101000000000000000010101";
                        f_reg(266) <= "00100011110111101111111111111111";
                        f_reg(267) <= "00100011111111111111111111111111";
                        f_reg(268) <= "00010111110111110000000001111101";
                        f_reg(269) <= "00011111111000001111111101001000";
                        f_reg(270) <= "00010000000000000000000100001000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "10001100000111010000011111001000";
                        f_reg(287) <= "00011111101000000000000000000011";
                        f_reg(288) <= "00100000000111010000000000111100";
                        f_reg(289) <= "00010000000000000000000000000010";
                        f_reg(290) <= "00100000000111010000000000000000";
                        f_reg(291) <= "00010100001011110000000001100110";
                        f_reg(292) <= "10101111101000010000011101010000";
                        f_reg(293) <= "10001100000111010000011111001000";
                        f_reg(294) <= "00011111101000000000000000000011";
                        f_reg(295) <= "00100000000111010000000000111100";
                        f_reg(296) <= "00010000000000000000000000000010";
                        f_reg(297) <= "00100000000111010000000000000000";
                        f_reg(298) <= "00010100010100000000000001011111";
                        f_reg(299) <= "10101111101000100000011101010100";
                        f_reg(300) <= "10001100000111010000011111001000";
                        f_reg(301) <= "00011111101000000000000000000011";
                        f_reg(302) <= "00100000000111010000000000111100";
                        f_reg(303) <= "00010000000000000000000000000010";
                        f_reg(304) <= "00100000000111010000000000000000";
                        f_reg(305) <= "00010100011100010000000001011000";
                        f_reg(306) <= "10101111101000110000011101011000";
                        f_reg(307) <= "10001100000111010000011111001000";
                        f_reg(308) <= "00011111101000000000000000000011";
                        f_reg(309) <= "00100000000111010000000000111100";
                        f_reg(310) <= "00010000000000000000000000000010";
                        f_reg(311) <= "00100000000111010000000000000000";
                        f_reg(312) <= "00010100100100100000000001010001";
                        f_reg(313) <= "10101111101001000000011101011100";
                        f_reg(314) <= "10001100000111010000011111001000";
                        f_reg(315) <= "00011111101000000000000000000011";
                        f_reg(316) <= "00100000000111010000000000111100";
                        f_reg(317) <= "00010000000000000000000000000010";
                        f_reg(318) <= "00100000000111010000000000000000";
                        f_reg(319) <= "00010100101100110000000001001010";
                        f_reg(320) <= "10101111101001010000011101100000";
                        f_reg(321) <= "10001100000111010000011111001000";
                        f_reg(322) <= "00011111101000000000000000000011";
                        f_reg(323) <= "00100000000111010000000000111100";
                        f_reg(324) <= "00010000000000000000000000000010";
                        f_reg(325) <= "00100000000111010000000000000000";
                        f_reg(326) <= "00010100110101000000000001000011";
                        f_reg(327) <= "10101111101001100000011101100100";
                        f_reg(328) <= "10001100000111010000011111001000";
                        f_reg(329) <= "00011111101000000000000000000011";
                        f_reg(330) <= "00100000000111010000000000111100";
                        f_reg(331) <= "00010000000000000000000000000010";
                        f_reg(332) <= "00100000000111010000000000000000";
                        f_reg(333) <= "00010100111101010000000000111100";
                        f_reg(334) <= "10101111101001110000011101101000";
                        f_reg(335) <= "10001100000111010000011111001000";
                        f_reg(336) <= "00011111101000000000000000000011";
                        f_reg(337) <= "00100000000111010000000000111100";
                        f_reg(338) <= "00010000000000000000000000000010";
                        f_reg(339) <= "00100000000111010000000000000000";
                        f_reg(340) <= "00010101000101100000000000110101";
                        f_reg(341) <= "10101111101010000000011101101100";
                        f_reg(342) <= "10001100000111010000011111001000";
                        f_reg(343) <= "00011111101000000000000000000011";
                        f_reg(344) <= "00100000000111010000000000111100";
                        f_reg(345) <= "00010000000000000000000000000010";
                        f_reg(346) <= "00100000000111010000000000000000";
                        f_reg(347) <= "00010101001101110000000000101110";
                        f_reg(348) <= "10101111101010010000011101110000";
                        f_reg(349) <= "10001100000111010000011111001000";
                        f_reg(350) <= "00011111101000000000000000000011";
                        f_reg(351) <= "00100000000111010000000000111100";
                        f_reg(352) <= "00010000000000000000000000000010";
                        f_reg(353) <= "00100000000111010000000000000000";
                        f_reg(354) <= "00010101010110000000000000100111";
                        f_reg(355) <= "10101111101010100000011101110100";
                        f_reg(356) <= "10001100000111010000011111001000";
                        f_reg(357) <= "00011111101000000000000000000011";
                        f_reg(358) <= "00100000000111010000000000111100";
                        f_reg(359) <= "00010000000000000000000000000010";
                        f_reg(360) <= "00100000000111010000000000000000";
                        f_reg(361) <= "00010101011110010000000000100000";
                        f_reg(362) <= "10101111101010110000011101111000";
                        f_reg(363) <= "10001100000111010000011111001000";
                        f_reg(364) <= "00011111101000000000000000000011";
                        f_reg(365) <= "00100000000111010000000000111100";
                        f_reg(366) <= "00010000000000000000000000000010";
                        f_reg(367) <= "00100000000111010000000000000000";
                        f_reg(368) <= "00010101100110100000000000011001";
                        f_reg(369) <= "10101111101011000000011101111100";
                        f_reg(370) <= "10001100000111010000011111001000";
                        f_reg(371) <= "00011111101000000000000000000011";
                        f_reg(372) <= "00100000000111010000000000111100";
                        f_reg(373) <= "00010000000000000000000000000010";
                        f_reg(374) <= "00100000000111010000000000000000";
                        f_reg(375) <= "00010101101110110000000000010010";
                        f_reg(376) <= "10101111101011010000011110000000";
                        f_reg(377) <= "10001100000111010000011111001000";
                        f_reg(378) <= "00011111101000000000000000000011";
                        f_reg(379) <= "00100000000111010000000000111100";
                        f_reg(380) <= "00010000000000000000000000000010";
                        f_reg(381) <= "00100000000111010000000000000000";
                        f_reg(382) <= "00010101110111000000000000001011";
                        f_reg(383) <= "10101111101011100000011110000100";
                        f_reg(384) <= "10001100000111010000011111001000";
                        f_reg(385) <= "00011111101000000000000000000011";
                        f_reg(386) <= "00100000000111010000000000111100";
                        f_reg(387) <= "00010000000000000000000000000010";
                        f_reg(388) <= "00100000000111010000000000000000";
                        f_reg(389) <= "00010111110111110000000000000100";
                        f_reg(390) <= "10101111101111100000011110001000";
                        f_reg(391) <= "10101100000111010000011111001000";
                        f_reg(392) <= "00010000000000001111111110000010";
                        f_reg(393) <= "10001100000111010000011111001000";
                        f_reg(394) <= "10001111101000010000011101010000";
                        f_reg(395) <= "10001100000111010000011111001000";
                        f_reg(396) <= "10001111101011110000011101010000";
                        f_reg(397) <= "00010100001011111111111111111100";
                        f_reg(398) <= "10001100000111010000011111001000";
                        f_reg(399) <= "10001111101000100000011101010100";
                        f_reg(400) <= "10001100000111010000011111001000";
                        f_reg(401) <= "10001111101100000000011101010100";
                        f_reg(402) <= "00010100010100001111111111111100";
                        f_reg(403) <= "10001100000111010000011111001000";
                        f_reg(404) <= "10001111101000110000011101011000";
                        f_reg(405) <= "10001100000111010000011111001000";
                        f_reg(406) <= "10001111101100010000011101011000";
                        f_reg(407) <= "00010100011100011111111111111100";
                        f_reg(408) <= "10001100000111010000011111001000";
                        f_reg(409) <= "10001111101001000000011101011100";
                        f_reg(410) <= "10001100000111010000011111001000";
                        f_reg(411) <= "10001111101100100000011101011100";
                        f_reg(412) <= "00010100100100101111111111111100";
                        f_reg(413) <= "10001100000111010000011111001000";
                        f_reg(414) <= "10001111101001010000011101100000";
                        f_reg(415) <= "10001100000111010000011111001000";
                        f_reg(416) <= "10001111101100110000011101100000";
                        f_reg(417) <= "00010100101100111111111111111100";
                        f_reg(418) <= "10001100000111010000011111001000";
                        f_reg(419) <= "10001111101001100000011101100100";
                        f_reg(420) <= "10001100000111010000011111001000";
                        f_reg(421) <= "10001111101101000000011101100100";
                        f_reg(422) <= "00010100110101001111111111111100";
                        f_reg(423) <= "10001100000111010000011111001000";
                        f_reg(424) <= "10001111101001110000011101101000";
                        f_reg(425) <= "10001100000111010000011111001000";
                        f_reg(426) <= "10001111101101010000011101101000";
                        f_reg(427) <= "00010100111101011111111111111100";
                        f_reg(428) <= "10001100000111010000011111001000";
                        f_reg(429) <= "10001111101010000000011101101100";
                        f_reg(430) <= "10001100000111010000011111001000";
                        f_reg(431) <= "10001111101101100000011101101100";
                        f_reg(432) <= "00010101000101101111111111111100";
                        f_reg(433) <= "10001100000111010000011111001000";
                        f_reg(434) <= "10001111101010010000011101110000";
                        f_reg(435) <= "10001100000111010000011111001000";
                        f_reg(436) <= "10001111101101110000011101110000";
                        f_reg(437) <= "00010101001101111111111111111100";
                        f_reg(438) <= "10001100000111010000011111001000";
                        f_reg(439) <= "10001111101010100000011101110100";
                        f_reg(440) <= "10001100000111010000011111001000";
                        f_reg(441) <= "10001111101110000000011101110100";
                        f_reg(442) <= "00010101010110001111111111111100";
                        f_reg(443) <= "10001100000111010000011111001000";
                        f_reg(444) <= "10001111101010110000011101111000";
                        f_reg(445) <= "10001100000111010000011111001000";
                        f_reg(446) <= "10001111101110010000011101111000";
                        f_reg(447) <= "00010101011110011111111111111100";
                        f_reg(448) <= "10001100000111010000011111001000";
                        f_reg(449) <= "10001111101011000000011101111100";
                        f_reg(450) <= "10001100000111010000011111001000";
                        f_reg(451) <= "10001111101110100000011101111100";
                        f_reg(452) <= "00010101100110101111111111111100";
                        f_reg(453) <= "10001100000111010000011111001000";
                        f_reg(454) <= "10001111101011010000011110000000";
                        f_reg(455) <= "10001100000111010000011111001000";
                        f_reg(456) <= "10001111101110110000011110000000";
                        f_reg(457) <= "00010101101110111111111111111100";
                        f_reg(458) <= "10001100000111010000011111001000";
                        f_reg(459) <= "10001111101011100000011110000100";
                        f_reg(460) <= "10001100000111010000011111001000";
                        f_reg(461) <= "10001111101111000000011110000100";
                        f_reg(462) <= "00010101110111001111111111111100";
                        f_reg(463) <= "10001100000111010000011111001000";
                        f_reg(464) <= "10001111101111100000011110001000";
                        f_reg(465) <= "10001100000111010000011111001000";
                        f_reg(466) <= "10001111101111110000011110001000";
                        f_reg(467) <= "00010111110111111111111111111100";
                        f_reg(468) <= "00010000000000001111111100110110";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000001111100111";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                     when others =>
                        -- Error if this occurs as there should never be a write to this address
                        f_DONE <= '1';
                        f_MEM_READY <= '0';
                        f_data <= B"00000000000000000000000000000000";
                        ff_MEM_READY <= '0';
                        f_read <= '0';
                        f_write <= '0';
                        f_sw_instr <= '0';
                        f_lw_instr <= '0';
                        f_br_instr <= '0';
                        f_last_address <= (others => '0');
                        f_next_address <= (others => '0');
                        f_sw_address <= (others => '0');
                        f_lw_address <= (others => '0');
                        f_branch_address <= (others => '0');
                        f_error_detected <= '0';
                        f_error_flag <= '0';
                        f_error <= (others => '0');
                        f_reg(1) <= "00111100000111110000001111100111";
                        f_reg(2) <= "00000000000111111111110000000010";
                        f_reg(3) <= "00111100000000011011010000101011";
                        f_reg(4) <= "00000000001000000001000000101011";
                        f_reg(5) <= "00111000010000111100011011001011";
                        f_reg(6) <= "00000000011000100010000000000100";
                        f_reg(7) <= "00000000001000110010100000101010";
                        f_reg(8) <= "00101100100001100111001010011100";
                        f_reg(9) <= "00101100110001111101001000000111";
                        f_reg(10) <= "00000000111001110100000000100110";
                        f_reg(11) <= "00110100101010010110110010111101";
                        f_reg(12) <= "00000000010001010101000000000110";
                        f_reg(13) <= "00000000000001110101110010000000";
                        f_reg(14) <= "10101100000000110000010000111000";
                        f_reg(15) <= "00000000010010010110000000100010";
                        f_reg(16) <= "00000000100000000110100000100101";
                        f_reg(17) <= "00110100000011100111011010100001";
                        f_reg(18) <= "00000001100011010111100000101010";
                        f_reg(19) <= "00000001000011111000000000000110";
                        f_reg(20) <= "00000000010011111000100000100110";
                        f_reg(21) <= "00111100000100100010010111000101";
                        f_reg(22) <= "00000000000001011001110101000000";
                        f_reg(23) <= "00000001101011101010000000101011";
                        f_reg(24) <= "00000000010000101010100000100011";
                        f_reg(25) <= "00000000011011100111000000000100";
                        f_reg(26) <= "00100100011101101001011111000111";
                        f_reg(27) <= "00000010110100001011100000000110";
                        f_reg(28) <= "00110010100110000111111001111001";
                        f_reg(29) <= "00000000100110001100100000100011";
                        f_reg(30) <= "10101100000100100000010000111100";
                        f_reg(31) <= "00000001001101011101000000000111";
                        f_reg(32) <= "00100111010110111101000101111101";
                        f_reg(33) <= "00000011000010101110000000100101";
                        f_reg(34) <= "00110100101111010110100111001000";
                        f_reg(35) <= "10101100000111000000010001000000";
                        f_reg(36) <= "00000010111001101111000000000110";
                        f_reg(37) <= "00000011010101100000100000100101";
                        f_reg(38) <= "10101100000111000000010001000100";
                        f_reg(39) <= "00110011110011001010100010100010";
                        f_reg(40) <= "00000001001111010100000000101010";
                        f_reg(41) <= "00000001100001000010000000100110";
                        f_reg(42) <= "00000001110110110111100000101010";
                        f_reg(43) <= "00000001011100010001000000100011";
                        f_reg(44) <= "00000000000011000001100101000010";
                        f_reg(45) <= "00000001000100111000000000100010";
                        f_reg(46) <= "00000000100001111010000000100110";
                        f_reg(47) <= "00000000010011011001000000100001";
                        f_reg(48) <= "00000000111000011010100000000100";
                        f_reg(49) <= "00101100011010100110000110110111";
                        f_reg(50) <= "00000010101110010010100000100111";
                        f_reg(51) <= "00000000000000000000000000000000";
                        f_reg(52) <= "00101110011001100101110000011101";
                        f_reg(53) <= "00000010010001011011100000000100";
                        f_reg(54) <= "00101011011110100111010011110100";
                        f_reg(55) <= "00000000000011111011001110000010";
                        f_reg(56) <= "00000000000000000000000000000000";
                        f_reg(57) <= "10101100000100110000010001001000";
                        f_reg(58) <= "00110011010111001111100100000000";
                        f_reg(59) <= "00000010111101000100100000100111";
                        f_reg(60) <= "00111100000111011011111101100111";
                        f_reg(61) <= "00000001010100000111000000000111";
                        f_reg(62) <= "00000001110001100101100000100100";
                        f_reg(63) <= "00000000000000000000000000000000";
                        f_reg(64) <= "10101100000010110000010001001100";
                        f_reg(65) <= "00000010110101101000100000100110";
                        f_reg(66) <= "10101100000111100000010001010000";
                        f_reg(67) <= "00000000000000000110011000000000";
                        f_reg(68) <= "00100111101010000010000000101001";
                        f_reg(69) <= "00000010001110000010000000100111";
                        f_reg(70) <= "00000001101010000001000000000110";
                        f_reg(71) <= "00000000000000000000000000000000";
                        f_reg(72) <= "00000001100111000000100000100110";
                        f_reg(73) <= "00000000010000010011100000000100";
                        f_reg(74) <= "00000000000000000000000000000000";
                        f_reg(75) <= "10101100000010010000010001010100";
                        f_reg(76) <= "10101100000001110000010001011000";
                        f_reg(77) <= "10101100000001000000010001011100";
                        f_reg(78) <= "00100011111111111111111111111111";
                        f_reg(79) <= "00011111111000001111111110110100";
                        f_reg(80) <= "00010000000000000000000111000110";
                        f_reg(81) <= "00111100000111100000001111100111";
                        f_reg(82) <= "00111100000111110000001111100111";
                        f_reg(83) <= "00000000000111101111010000000010";
                        f_reg(84) <= "00000000000111111111110000000010";
                        f_reg(85) <= "00111100000000011011010000101011";
                        f_reg(86) <= "00111100000011111011010000101011";
                        f_reg(87) <= "00000000001000000001000000101011";
                        f_reg(88) <= "00000001111000001000000000101011";
                        f_reg(89) <= "00111000010000111100011011001011";
                        f_reg(90) <= "00111010000100011100011011001011";
                        f_reg(91) <= "00000000011000100010000000000100";
                        f_reg(92) <= "00000010001100001001000000000100";
                        f_reg(93) <= "00000000001000110010100000101010";
                        f_reg(94) <= "00000001111100011001100000101010";
                        f_reg(95) <= "00101100100001100111001010011100";
                        f_reg(96) <= "00101110010101000111001010011100";
                        f_reg(97) <= "00101100110001111101001000000111";
                        f_reg(98) <= "00101110100101011101001000000111";
                        f_reg(99) <= "00000000111001110100000000100110";
                        f_reg(100) <= "00000010101101011011000000100110";
                        f_reg(101) <= "00110100101010010110110010111101";
                        f_reg(102) <= "00110110011101110110110010111101";
                        f_reg(103) <= "00000000010001010101000000000110";
                        f_reg(104) <= "00000010000100111100000000000110";
                        f_reg(105) <= "00000000000001110101110010000000";
                        f_reg(106) <= "00000000000101011100110010000000";
                        f_reg(107) <= "00010100011100010000000100011110";
                        f_reg(108) <= "10101100000000110000010000111000";
                        f_reg(109) <= "00000000010010010110000000100010";
                        f_reg(110) <= "00000010000101111101000000100010";
                        f_reg(111) <= "00000000100000000110100000100101";
                        f_reg(112) <= "00000010010000001101100000100101";
                        f_reg(113) <= "00110100000011100111011010100001";
                        f_reg(114) <= "00110100000111000111011010100001";
                        f_reg(115) <= "00000001100011010000100000101010";
                        f_reg(116) <= "00000011010110110111100000101010";
                        f_reg(117) <= "00000001000000010110000000000110";
                        f_reg(118) <= "00000010110011111101000000000110";
                        f_reg(119) <= "00000000010000010100000000100110";
                        f_reg(120) <= "00000010000011111011000000100110";
                        f_reg(121) <= "00111100000000010010010111000101";
                        f_reg(122) <= "00111100000011110010010111000101";
                        f_reg(123) <= "00010101101110110000000100001110";
                        f_reg(124) <= "10101100000011010000010001100000";
                        f_reg(125) <= "00000000000001010110110101000000";
                        f_reg(126) <= "00000000000100111101110101000000";
                        f_reg(127) <= "00010101101110110000000100001010";
                        f_reg(128) <= "10101100000011010000010001100100";
                        f_reg(129) <= "10001100000011010000010001100000";
                        f_reg(130) <= "10001100000110110000010001100000";
                        f_reg(131) <= "00010101101110111111111111111110";
                        f_reg(132) <= "00010100111101010000000100000101";
                        f_reg(133) <= "10101100000001110000010001101000";
                        f_reg(134) <= "00000001101011100011100000101011";
                        f_reg(135) <= "00000011011111001010100000101011";
                        f_reg(136) <= "00010101101110110000000100000001";
                        f_reg(137) <= "10101100000011010000010001101100";
                        f_reg(138) <= "00000000010000100110100000100011";
                        f_reg(139) <= "00000010000100001101100000100011";
                        f_reg(140) <= "00000000011011100111000000000100";
                        f_reg(141) <= "00000010001111001110000000000100";
                        f_reg(142) <= "00100100011000101001011111000111";
                        f_reg(143) <= "00100110001100001001011111000111";
                        f_reg(144) <= "00000000010011000001100000000110";
                        f_reg(145) <= "00000010000110101000100000000110";
                        f_reg(146) <= "00110000111011000111111001111001";
                        f_reg(147) <= "00110010101110100111111001111001";
                        f_reg(148) <= "00000000100011000011100000100011";
                        f_reg(149) <= "00000010010110101010100000100011";
                        f_reg(150) <= "00010100001011110000000011110011";
                        f_reg(151) <= "10101100000000010000010000111100";
                        f_reg(152) <= "00000001001011010000100000000111";
                        f_reg(153) <= "00000010111110110111100000000111";
                        f_reg(154) <= "00100100001011011101000101111101";
                        f_reg(155) <= "00100101111110111101000101111101";
                        f_reg(156) <= "00010101101110110000000011101101";
                        f_reg(157) <= "10101100000011010000010001110000";
                        f_reg(158) <= "00000001100010100110100000100101";
                        f_reg(159) <= "00000011010110001101100000100101";
                        f_reg(160) <= "00110100101010100110100111001000";
                        f_reg(161) <= "00110110011110000110100111001000";
                        f_reg(162) <= "00010101101110110000000011100111";
                        f_reg(163) <= "10101100000011010000010001000000";
                        f_reg(164) <= "00000000011001100010100000000110";
                        f_reg(165) <= "00000010001101001001100000000110";
                        f_reg(166) <= "00000000001000100011000000100101";
                        f_reg(167) <= "00000001111100001010000000100101";
                        f_reg(168) <= "00010101101110110000000011100001";
                        f_reg(169) <= "10101100000011010000010001000100";
                        f_reg(170) <= "00110000101000111010100010100010";
                        f_reg(171) <= "00110010011100011010100010100010";
                        f_reg(172) <= "00000001001010100000100000101010";
                        f_reg(173) <= "00000010111110000111100000101010";
                        f_reg(174) <= "00000000011001000010000000100110";
                        f_reg(175) <= "00000010001100101001000000100110";
                        f_reg(176) <= "10001100000000100000010001110000";
                        f_reg(177) <= "10001100000100000000010001110000";
                        f_reg(178) <= "00010100010100001111111111111110";
                        f_reg(179) <= "00000001110000100110100000101010";
                        f_reg(180) <= "00000011100100001101100000101010";
                        f_reg(181) <= "00000001011010000100100000100011";
                        f_reg(182) <= "00000011001101101011100000100011";
                        f_reg(183) <= "00000000000000110101000101000010";
                        f_reg(184) <= "00000000000100011100000101000010";
                        f_reg(185) <= "10001100000011100000010001100100";
                        f_reg(186) <= "10001100000111000000010001100100";
                        f_reg(187) <= "00010101110111001111111111111110";
                        f_reg(188) <= "00000000001011100101100000100010";
                        f_reg(189) <= "00000001111111001100100000100010";
                        f_reg(190) <= "10001100000010000000010001101000";
                        f_reg(191) <= "10001100000101100000010001101000";
                        f_reg(192) <= "00010101000101101111111111111110";
                        f_reg(193) <= "00000000100010000001100000100110";
                        f_reg(194) <= "00000010010101101000100000100110";
                        f_reg(195) <= "10001100000000010000010001101100";
                        f_reg(196) <= "10001100000011110000010001101100";
                        f_reg(197) <= "00010100001011111111111111111110";
                        f_reg(198) <= "00000001001000010010000000100001";
                        f_reg(199) <= "00000010111011111001000000100001";
                        f_reg(200) <= "00000001000001100100100000000100";
                        f_reg(201) <= "00000010110101001011100000000100";
                        f_reg(202) <= "00101101010001100110000110110111";
                        f_reg(203) <= "00101111000101000110000110110111";
                        f_reg(204) <= "00000001001001110100000000100111";
                        f_reg(205) <= "00000010111101011011000000100111";
                        f_reg(206) <= "00000000000000000000000000000000";
                        f_reg(207) <= "00000000000000000000000000000000";
                        f_reg(208) <= "00101101110010100101110000011101";
                        f_reg(209) <= "00101111100110000101110000011101";
                        f_reg(210) <= "00000000100010000100100000000100";
                        f_reg(211) <= "00000010010101101011100000000100";
                        f_reg(212) <= "00101000010001110111010011110100";
                        f_reg(213) <= "00101010000101010111010011110100";
                        f_reg(214) <= "00000000000011010100001110000010";
                        f_reg(215) <= "00000000000110111011001110000010";
                        f_reg(216) <= "00000000000000000000000000000000";
                        f_reg(217) <= "00000000000000000000000000000000";
                        f_reg(218) <= "00010101110111000000000010101111";
                        f_reg(219) <= "10101100000011100000010001001000";
                        f_reg(220) <= "00110000111001001111100100000000";
                        f_reg(221) <= "00110010101100101111100100000000";
                        f_reg(222) <= "00000001001000110001000000100111";
                        f_reg(223) <= "00000010111100011000000000100111";
                        f_reg(224) <= "00111100000011011011111101100111";
                        f_reg(225) <= "00111100000110111011111101100111";
                        f_reg(226) <= "00000000110010110111000000000111";
                        f_reg(227) <= "00000010100110011110000000000111";
                        f_reg(228) <= "00000001110010100011100000100100";
                        f_reg(229) <= "00000011100110001010100000100100";
                        f_reg(230) <= "00000000000000000000000000000000";
                        f_reg(231) <= "00000000000000000000000000000000";
                        f_reg(232) <= "00010100111101010000000010100001";
                        f_reg(233) <= "10101100000001110000010001001100";
                        f_reg(234) <= "00000001000010000100100000100110";
                        f_reg(235) <= "00000010110101101011100000100110";
                        f_reg(236) <= "00010100101100110000000010011101";
                        f_reg(237) <= "10101100000001010000010001010000";
                        f_reg(238) <= "00000000000000000001111000000000";
                        f_reg(239) <= "00000000000000001000111000000000";
                        f_reg(240) <= "00100101101010110010000000101001";
                        f_reg(241) <= "00100111011110010010000000101001";
                        f_reg(242) <= "00000001001011000011000000100111";
                        f_reg(243) <= "00000010111110101010000000100111";
                        f_reg(244) <= "00000000001010110111000000000110";
                        f_reg(245) <= "00000001111110011110000000000110";
                        f_reg(246) <= "00000000000000000000000000000000";
                        f_reg(247) <= "00000000000000000000000000000000";
                        f_reg(248) <= "00000000011001000101000000100110";
                        f_reg(249) <= "00000010001100101100000000100110";
                        f_reg(250) <= "00000001110010100011100000000100";
                        f_reg(251) <= "00000011100110001010100000000100";
                        f_reg(252) <= "00000000000000000000000000000000";
                        f_reg(253) <= "00000000000000000000000000000000";
                        f_reg(254) <= "00010100010100000000000010001011";
                        f_reg(255) <= "10101100000000100000010001010100";
                        f_reg(256) <= "00010100111101010000000010001001";
                        f_reg(257) <= "10101100000001110000010001011000";
                        f_reg(258) <= "00010100110101000000000010000111";
                        f_reg(259) <= "10101100000001100000010001011100";
                        f_reg(260) <= "00100011110111011111111100000110";
                        f_reg(261) <= "00010011101000000000000000011001";
                        f_reg(262) <= "00100011110111011111111000001100";
                        f_reg(263) <= "00010011101000000000000000010111";
                        f_reg(264) <= "00100011110111011111110100010010";
                        f_reg(265) <= "00010011101000000000000000010101";
                        f_reg(266) <= "00100011110111101111111111111111";
                        f_reg(267) <= "00100011111111111111111111111111";
                        f_reg(268) <= "00010111110111110000000001111101";
                        f_reg(269) <= "00011111111000001111111101001000";
                        f_reg(270) <= "00010000000000000000000100001000";
                        f_reg(271) <= "00000000000000000000000000000000";
                        f_reg(272) <= "00000000000000000000000000000000";
                        f_reg(273) <= "00000000000000000000000000000000";
                        f_reg(274) <= "00000000000000000000000000000000";
                        f_reg(275) <= "00000000000000000000000000000000";
                        f_reg(276) <= "00000000000000000000000000000000";
                        f_reg(277) <= "00000000000000000000000000000000";
                        f_reg(278) <= "00000000000000000000000000000000";
                        f_reg(279) <= "00000000000000000000000000000000";
                        f_reg(280) <= "00000000000000000000000000000000";
                        f_reg(281) <= "00000000000000000000000000000000";
                        f_reg(282) <= "00000000000000000000000000000000";
                        f_reg(283) <= "00000000000000000000000000000000";
                        f_reg(284) <= "00000000000000000000000000000000";
                        f_reg(285) <= "00000000000000000000000000000000";
                        f_reg(286) <= "10001100000111010000011111001000";
                        f_reg(287) <= "00011111101000000000000000000011";
                        f_reg(288) <= "00100000000111010000000000111100";
                        f_reg(289) <= "00010000000000000000000000000010";
                        f_reg(290) <= "00100000000111010000000000000000";
                        f_reg(291) <= "00010100001011110000000001100110";
                        f_reg(292) <= "10101111101000010000011101010000";
                        f_reg(293) <= "10001100000111010000011111001000";
                        f_reg(294) <= "00011111101000000000000000000011";
                        f_reg(295) <= "00100000000111010000000000111100";
                        f_reg(296) <= "00010000000000000000000000000010";
                        f_reg(297) <= "00100000000111010000000000000000";
                        f_reg(298) <= "00010100010100000000000001011111";
                        f_reg(299) <= "10101111101000100000011101010100";
                        f_reg(300) <= "10001100000111010000011111001000";
                        f_reg(301) <= "00011111101000000000000000000011";
                        f_reg(302) <= "00100000000111010000000000111100";
                        f_reg(303) <= "00010000000000000000000000000010";
                        f_reg(304) <= "00100000000111010000000000000000";
                        f_reg(305) <= "00010100011100010000000001011000";
                        f_reg(306) <= "10101111101000110000011101011000";
                        f_reg(307) <= "10001100000111010000011111001000";
                        f_reg(308) <= "00011111101000000000000000000011";
                        f_reg(309) <= "00100000000111010000000000111100";
                        f_reg(310) <= "00010000000000000000000000000010";
                        f_reg(311) <= "00100000000111010000000000000000";
                        f_reg(312) <= "00010100100100100000000001010001";
                        f_reg(313) <= "10101111101001000000011101011100";
                        f_reg(314) <= "10001100000111010000011111001000";
                        f_reg(315) <= "00011111101000000000000000000011";
                        f_reg(316) <= "00100000000111010000000000111100";
                        f_reg(317) <= "00010000000000000000000000000010";
                        f_reg(318) <= "00100000000111010000000000000000";
                        f_reg(319) <= "00010100101100110000000001001010";
                        f_reg(320) <= "10101111101001010000011101100000";
                        f_reg(321) <= "10001100000111010000011111001000";
                        f_reg(322) <= "00011111101000000000000000000011";
                        f_reg(323) <= "00100000000111010000000000111100";
                        f_reg(324) <= "00010000000000000000000000000010";
                        f_reg(325) <= "00100000000111010000000000000000";
                        f_reg(326) <= "00010100110101000000000001000011";
                        f_reg(327) <= "10101111101001100000011101100100";
                        f_reg(328) <= "10001100000111010000011111001000";
                        f_reg(329) <= "00011111101000000000000000000011";
                        f_reg(330) <= "00100000000111010000000000111100";
                        f_reg(331) <= "00010000000000000000000000000010";
                        f_reg(332) <= "00100000000111010000000000000000";
                        f_reg(333) <= "00010100111101010000000000111100";
                        f_reg(334) <= "10101111101001110000011101101000";
                        f_reg(335) <= "10001100000111010000011111001000";
                        f_reg(336) <= "00011111101000000000000000000011";
                        f_reg(337) <= "00100000000111010000000000111100";
                        f_reg(338) <= "00010000000000000000000000000010";
                        f_reg(339) <= "00100000000111010000000000000000";
                        f_reg(340) <= "00010101000101100000000000110101";
                        f_reg(341) <= "10101111101010000000011101101100";
                        f_reg(342) <= "10001100000111010000011111001000";
                        f_reg(343) <= "00011111101000000000000000000011";
                        f_reg(344) <= "00100000000111010000000000111100";
                        f_reg(345) <= "00010000000000000000000000000010";
                        f_reg(346) <= "00100000000111010000000000000000";
                        f_reg(347) <= "00010101001101110000000000101110";
                        f_reg(348) <= "10101111101010010000011101110000";
                        f_reg(349) <= "10001100000111010000011111001000";
                        f_reg(350) <= "00011111101000000000000000000011";
                        f_reg(351) <= "00100000000111010000000000111100";
                        f_reg(352) <= "00010000000000000000000000000010";
                        f_reg(353) <= "00100000000111010000000000000000";
                        f_reg(354) <= "00010101010110000000000000100111";
                        f_reg(355) <= "10101111101010100000011101110100";
                        f_reg(356) <= "10001100000111010000011111001000";
                        f_reg(357) <= "00011111101000000000000000000011";
                        f_reg(358) <= "00100000000111010000000000111100";
                        f_reg(359) <= "00010000000000000000000000000010";
                        f_reg(360) <= "00100000000111010000000000000000";
                        f_reg(361) <= "00010101011110010000000000100000";
                        f_reg(362) <= "10101111101010110000011101111000";
                        f_reg(363) <= "10001100000111010000011111001000";
                        f_reg(364) <= "00011111101000000000000000000011";
                        f_reg(365) <= "00100000000111010000000000111100";
                        f_reg(366) <= "00010000000000000000000000000010";
                        f_reg(367) <= "00100000000111010000000000000000";
                        f_reg(368) <= "00010101100110100000000000011001";
                        f_reg(369) <= "10101111101011000000011101111100";
                        f_reg(370) <= "10001100000111010000011111001000";
                        f_reg(371) <= "00011111101000000000000000000011";
                        f_reg(372) <= "00100000000111010000000000111100";
                        f_reg(373) <= "00010000000000000000000000000010";
                        f_reg(374) <= "00100000000111010000000000000000";
                        f_reg(375) <= "00010101101110110000000000010010";
                        f_reg(376) <= "10101111101011010000011110000000";
                        f_reg(377) <= "10001100000111010000011111001000";
                        f_reg(378) <= "00011111101000000000000000000011";
                        f_reg(379) <= "00100000000111010000000000111100";
                        f_reg(380) <= "00010000000000000000000000000010";
                        f_reg(381) <= "00100000000111010000000000000000";
                        f_reg(382) <= "00010101110111000000000000001011";
                        f_reg(383) <= "10101111101011100000011110000100";
                        f_reg(384) <= "10001100000111010000011111001000";
                        f_reg(385) <= "00011111101000000000000000000011";
                        f_reg(386) <= "00100000000111010000000000111100";
                        f_reg(387) <= "00010000000000000000000000000010";
                        f_reg(388) <= "00100000000111010000000000000000";
                        f_reg(389) <= "00010111110111110000000000000100";
                        f_reg(390) <= "10101111101111100000011110001000";
                        f_reg(391) <= "10101100000111010000011111001000";
                        f_reg(392) <= "00010000000000001111111110000010";
                        f_reg(393) <= "10001100000111010000011111001000";
                        f_reg(394) <= "10001111101000010000011101010000";
                        f_reg(395) <= "10001100000111010000011111001000";
                        f_reg(396) <= "10001111101011110000011101010000";
                        f_reg(397) <= "00010100001011111111111111111100";
                        f_reg(398) <= "10001100000111010000011111001000";
                        f_reg(399) <= "10001111101000100000011101010100";
                        f_reg(400) <= "10001100000111010000011111001000";
                        f_reg(401) <= "10001111101100000000011101010100";
                        f_reg(402) <= "00010100010100001111111111111100";
                        f_reg(403) <= "10001100000111010000011111001000";
                        f_reg(404) <= "10001111101000110000011101011000";
                        f_reg(405) <= "10001100000111010000011111001000";
                        f_reg(406) <= "10001111101100010000011101011000";
                        f_reg(407) <= "00010100011100011111111111111100";
                        f_reg(408) <= "10001100000111010000011111001000";
                        f_reg(409) <= "10001111101001000000011101011100";
                        f_reg(410) <= "10001100000111010000011111001000";
                        f_reg(411) <= "10001111101100100000011101011100";
                        f_reg(412) <= "00010100100100101111111111111100";
                        f_reg(413) <= "10001100000111010000011111001000";
                        f_reg(414) <= "10001111101001010000011101100000";
                        f_reg(415) <= "10001100000111010000011111001000";
                        f_reg(416) <= "10001111101100110000011101100000";
                        f_reg(417) <= "00010100101100111111111111111100";
                        f_reg(418) <= "10001100000111010000011111001000";
                        f_reg(419) <= "10001111101001100000011101100100";
                        f_reg(420) <= "10001100000111010000011111001000";
                        f_reg(421) <= "10001111101101000000011101100100";
                        f_reg(422) <= "00010100110101001111111111111100";
                        f_reg(423) <= "10001100000111010000011111001000";
                        f_reg(424) <= "10001111101001110000011101101000";
                        f_reg(425) <= "10001100000111010000011111001000";
                        f_reg(426) <= "10001111101101010000011101101000";
                        f_reg(427) <= "00010100111101011111111111111100";
                        f_reg(428) <= "10001100000111010000011111001000";
                        f_reg(429) <= "10001111101010000000011101101100";
                        f_reg(430) <= "10001100000111010000011111001000";
                        f_reg(431) <= "10001111101101100000011101101100";
                        f_reg(432) <= "00010101000101101111111111111100";
                        f_reg(433) <= "10001100000111010000011111001000";
                        f_reg(434) <= "10001111101010010000011101110000";
                        f_reg(435) <= "10001100000111010000011111001000";
                        f_reg(436) <= "10001111101101110000011101110000";
                        f_reg(437) <= "00010101001101111111111111111100";
                        f_reg(438) <= "10001100000111010000011111001000";
                        f_reg(439) <= "10001111101010100000011101110100";
                        f_reg(440) <= "10001100000111010000011111001000";
                        f_reg(441) <= "10001111101110000000011101110100";
                        f_reg(442) <= "00010101010110001111111111111100";
                        f_reg(443) <= "10001100000111010000011111001000";
                        f_reg(444) <= "10001111101010110000011101111000";
                        f_reg(445) <= "10001100000111010000011111001000";
                        f_reg(446) <= "10001111101110010000011101111000";
                        f_reg(447) <= "00010101011110011111111111111100";
                        f_reg(448) <= "10001100000111010000011111001000";
                        f_reg(449) <= "10001111101011000000011101111100";
                        f_reg(450) <= "10001100000111010000011111001000";
                        f_reg(451) <= "10001111101110100000011101111100";
                        f_reg(452) <= "00010101100110101111111111111100";
                        f_reg(453) <= "10001100000111010000011111001000";
                        f_reg(454) <= "10001111101011010000011110000000";
                        f_reg(455) <= "10001100000111010000011111001000";
                        f_reg(456) <= "10001111101110110000011110000000";
                        f_reg(457) <= "00010101101110111111111111111100";
                        f_reg(458) <= "10001100000111010000011111001000";
                        f_reg(459) <= "10001111101011100000011110000100";
                        f_reg(460) <= "10001100000111010000011111001000";
                        f_reg(461) <= "10001111101111000000011110000100";
                        f_reg(462) <= "00010101110111001111111111111100";
                        f_reg(463) <= "10001100000111010000011111001000";
                        f_reg(464) <= "10001111101111100000011110001000";
                        f_reg(465) <= "10001100000111010000011111001000";
                        f_reg(466) <= "10001111101111110000011110001000";
                        f_reg(467) <= "00010111110111111111111111111100";
                        f_reg(468) <= "00010000000000001111111100110110";
                        f_reg(469) <= "00000000000000000000000000000000";
                        f_reg(470) <= "00000000000000000000000000000000";
                        f_reg(471) <= "00000000000000000000000000000000";
                        f_reg(472) <= "00000000000000000000000000000000";
                        f_reg(473) <= "00000000000000000000000000000000";
                        f_reg(474) <= "00000000000000000000000000000000";
                        f_reg(475) <= "00000000000000000000000000000000";
                        f_reg(476) <= "00000000000000000000000000000000";
                        f_reg(477) <= "00000000000000000000000000000000";
                        f_reg(478) <= "00000000000000000000000000000000";
                        f_reg(479) <= "00000000000000000000000000000000";
                        f_reg(480) <= "00000000000000000000000000000000";
                        f_reg(481) <= "00000000000000000000000000000000";
                        f_reg(482) <= "00000000000000000000000000000000";
                        f_reg(483) <= "00000000000000000000000000000000";
                        f_reg(484) <= "00000000000000000000000000000000";
                        f_reg(485) <= "00000000000000000000000000000000";
                        f_reg(486) <= "00000000000000000000000000000000";
                        f_reg(487) <= "00000000000000000000000000000000";
                        f_reg(488) <= "00000000000000000000000000000000";
                        f_reg(489) <= "00000000000000000000000000000000";
                        f_reg(490) <= "00000000000000000000000000000000";
                        f_reg(491) <= "00000000000000000000000000000000";
                        f_reg(492) <= "00000000000000000000000000000000";
                        f_reg(493) <= "00000000000000000000000000000000";
                        f_reg(494) <= "00000000000000000000000000000000";
                        f_reg(495) <= "00000000000000000000000000000000";
                        f_reg(496) <= "00000000000000000000000000000000";
                        f_reg(497) <= "00000000000000000000000000000000";
                        f_reg(498) <= "00000000000000000000000000000000";
                        f_reg(499) <= "00000000000000000000001111100111";
                        f_reg(500) <= "00000000000000000000000000000000";
                        f_reg(501) <= "00000000000000000000000000000000";
                        f_reg(502) <= "00000000000000000000000000000000";
                        f_reg(503) <= "00000000000000000000000000000000";
                        f_reg(504) <= "00000000000000000000000000000000";
                        f_reg(505) <= "00000000000000000000000000000000";
                        f_reg(506) <= "00000000000000000000000000000000";
                        f_reg(507) <= "00000000000000000000000000000000";
                        f_reg(508) <= "00000000000000000000000000000000";
                        f_reg(509) <= "00000000000000000000000000000000";
                        f_reg(510) <= "00000000000000000000000000000000";
                        f_reg(511) <= "00000000000000000000000000000000";
                        f_reg(512) <= "00000000000000000000000000000000";
                        f_reg(513) <= "00000000000000000000000000000000";
                        f_reg(514) <= "00000000000000000000000000000000";
                        f_reg(515) <= "00000000000000000000000000000000";
                        f_reg(516) <= "00000000000000000000000000000000";
                        f_reg(517) <= "00000000000000000000000000000000";
                        f_reg(518) <= "00000000000000000000000000000000";
                        f_reg(519) <= "00000000000000000000000000000000";
                        f_reg(520) <= "00000000000000000000000000000000";
                        f_reg(521) <= "00000000000000000000000000000000";
                        f_reg(522) <= "00000000000000000000000000000000";
                        f_reg(523) <= "00000000000000000000000000000000";
                        f_reg(524) <= "00000000000000000000000000000000";
                        f_reg(525) <= "00000000000000000000000000000000";
                        f_reg(526) <= "00000000000000000000000000000000";
                        f_reg(527) <= "00000000000000000000000000000000";
                        f_reg(528) <= "00000000000000000000000000000000";
                        f_reg(529) <= "00000000000000000000000000000000";
                        f_reg(530) <= "00000000000000000000000000000000";
                        f_reg(531) <= "00000000000000000000000000000000";
                        f_reg(532) <= "00000000000000000000000000000000";
                        f_reg(533) <= "00000000000000000000000000000000";
                  end case;
               -- Data request already received.  Conitnue providing same outputs
               else
                  f_MEM_READY <= f_MEM_READY;
               end if;

            -- Not attempting to read from or write to memory
            else
               f_read <= '0';
               f_write <= '0';
               f_MEM_READY <= '0';
            end if;
         else
            f_DONE <= '0';
         end if;
      end if;
   end process;
end a_Test79_Reg_COMBINED;
